/*
Signal Generator - Creates a sine wave that has the supplied input frequency.
	Operates from 100Hz to 8000Hz.  
	
	outputSample is the current sine amplitude.
	
	
	This is a bit hardcoded to 128 total samples at a 32000 clock but can be changed by modifying some of the constants.
*/

module SignalGenerator_Bee  ( 
		input logic CLK_32KHz,
		input logic reset_n,
		input logic[13:0] inputFrequency,
		input logic [7:0] inputAmplitude, //Can give it a constant amplitude as well
		input logic [7:0] inputOffset, //Offset starting value
		output logic[7 : 0] outputSample,
		output logic indexZero
		);
		

	//Will count up to 320000.
	reg [20 : 0] counter ; //16 bits max value is 64k ~
	reg [7:0] smoothAmplitude;
	reg [10:0] smoothAmpCounter;

	always_ff @(posedge CLK_32KHz, negedge reset_n) begin
		if (reset_n == 1'b0)begin
			counter <= inputOffset * 125;
			smoothAmpCounter <= 0;
			smoothAmplitude <= 0;
		end
		else begin
			//If counter reaches top of index, it gets reduced by 32000 but keeps whatever it overshot by.  
			if (counter == (16'd66996)) begin  counter <= 66996; end
			//if (counter >= (16'd66996)) begin  counter <= counter - (16'd66996 ) + inputFrequency; end
			//inputFrequency holds 14 bits, so we need 2 extra in front.
			else begin counter <= counter + (inputFrequency);end//{ 2'b0, inputFrequency }; end

			if (smoothAmpCounter == 100)  begin
				smoothAmpCounter <= 0;
				if (smoothAmplitude < inputAmplitude) begin smoothAmplitude <= smoothAmplitude + 1; end
				else if (smoothAmplitude > inputAmplitude) begin smoothAmplitude <= smoothAmplitude - 1; end
			end 
			else begin
				smoothAmpCounter <= smoothAmpCounter + 1;
			end
		end
	end

	wire [20:0] trueCounter ;

	assign trueCounter = ( ( (counter/16) % 16'd16749) ) ;   // 0.trueCounter == 1/252 
	assign outputSample =  SignalMultiply255(soundFileAmplitudes[trueCounter],smoothAmplitude );   //Combine amplitude with input.  
	assign indexZero = (trueCounter == 0) ? 1'b1 : 1'b0;

	//Combines tow signals into 1
	function automatic  [7:0] SignalMultiply255 (input [7:0] a, input [7:0] b);
		return  ( (a * b + 127) * 1/255);
	endfunction		

	//--------------------------------------------
	//  [Amount of bits -1] Name [AmountOfSamples]//COPY PASTE FROM FILE STARTING ON THIS LINE DOWNWARD. INCLUDE ENDMODULE
bit [16749:0][7:0] soundFileAmplitudes;

//-=-=-=-=-SONG DATA-=-=-=-=- 
   assign soundFileAmplitudes [0] = 8'd123;
   assign soundFileAmplitudes [1] = 8'd134;
   assign soundFileAmplitudes [2] = 8'd151;
   assign soundFileAmplitudes [3] = 8'd155;
   assign soundFileAmplitudes [4] = 8'd144;
   assign soundFileAmplitudes [5] = 8'd128;
   assign soundFileAmplitudes [6] = 8'd117;
   assign soundFileAmplitudes [7] = 8'd105;
   assign soundFileAmplitudes [8] = 8'd106;
   assign soundFileAmplitudes [9] = 8'd113;
   assign soundFileAmplitudes [10] = 8'd116;
   assign soundFileAmplitudes [11] = 8'd125;
   assign soundFileAmplitudes [12] = 8'd128;
   assign soundFileAmplitudes [13] = 8'd118;
   assign soundFileAmplitudes [14] = 8'd120;
   assign soundFileAmplitudes [15] = 8'd118;
   assign soundFileAmplitudes [16] = 8'd122;
   assign soundFileAmplitudes [17] = 8'd137;
   assign soundFileAmplitudes [18] = 8'd146;
   assign soundFileAmplitudes [19] = 8'd152;
   assign soundFileAmplitudes [20] = 8'd147;
   assign soundFileAmplitudes [21] = 8'd141;
   assign soundFileAmplitudes [22] = 8'd144;
   assign soundFileAmplitudes [23] = 8'd136;
   assign soundFileAmplitudes [24] = 8'd125;
   assign soundFileAmplitudes [25] = 8'd123;
   assign soundFileAmplitudes [26] = 8'd120;
   assign soundFileAmplitudes [27] = 8'd114;
   assign soundFileAmplitudes [28] = 8'd96;
   assign soundFileAmplitudes [29] = 8'd75;
   assign soundFileAmplitudes [30] = 8'd90;
   assign soundFileAmplitudes [31] = 8'd115;
   assign soundFileAmplitudes [32] = 8'd126;
   assign soundFileAmplitudes [33] = 8'd132;
   assign soundFileAmplitudes [34] = 8'd131;
   assign soundFileAmplitudes [35] = 8'd133;
   assign soundFileAmplitudes [36] = 8'd146;
   assign soundFileAmplitudes [37] = 8'd163;
   assign soundFileAmplitudes [38] = 8'd154;
   assign soundFileAmplitudes [39] = 8'd138;
   assign soundFileAmplitudes [40] = 8'd137;
   assign soundFileAmplitudes [41] = 8'd127;
   assign soundFileAmplitudes [42] = 8'd112;
   assign soundFileAmplitudes [43] = 8'd107;
   assign soundFileAmplitudes [44] = 8'd104;
   assign soundFileAmplitudes [45] = 8'd106;
   assign soundFileAmplitudes [46] = 8'd114;
   assign soundFileAmplitudes [47] = 8'd121;
   assign soundFileAmplitudes [48] = 8'd128;
   assign soundFileAmplitudes [49] = 8'd133;
   assign soundFileAmplitudes [50] = 8'd131;
   assign soundFileAmplitudes [51] = 8'd134;
   assign soundFileAmplitudes [52] = 8'd143;
   assign soundFileAmplitudes [53] = 8'd157;
   assign soundFileAmplitudes [54] = 8'd160;
   assign soundFileAmplitudes [55] = 8'd140;
   assign soundFileAmplitudes [56] = 8'd141;
   assign soundFileAmplitudes [57] = 8'd139;
   assign soundFileAmplitudes [58] = 8'd122;
   assign soundFileAmplitudes [59] = 8'd111;
   assign soundFileAmplitudes [60] = 8'd105;
   assign soundFileAmplitudes [61] = 8'd103;
   assign soundFileAmplitudes [62] = 8'd94;
   assign soundFileAmplitudes [63] = 8'd87;
   assign soundFileAmplitudes [64] = 8'd90;
   assign soundFileAmplitudes [65] = 8'd108;
   assign soundFileAmplitudes [66] = 8'd129;
   assign soundFileAmplitudes [67] = 8'd137;
   assign soundFileAmplitudes [68] = 8'd135;
   assign soundFileAmplitudes [69] = 8'd127;
   assign soundFileAmplitudes [70] = 8'd138;
   assign soundFileAmplitudes [71] = 8'd155;
   assign soundFileAmplitudes [72] = 8'd155;
   assign soundFileAmplitudes [73] = 8'd142;
   assign soundFileAmplitudes [74] = 8'd128;
   assign soundFileAmplitudes [75] = 8'd126;
   assign soundFileAmplitudes [76] = 8'd103;
   assign soundFileAmplitudes [77] = 8'd112;
   assign soundFileAmplitudes [78] = 8'd123;
   assign soundFileAmplitudes [79] = 8'd130;
   assign soundFileAmplitudes [80] = 8'd138;
   assign soundFileAmplitudes [81] = 8'd126;
   assign soundFileAmplitudes [82] = 8'd125;
   assign soundFileAmplitudes [83] = 8'd130;
   assign soundFileAmplitudes [84] = 8'd130;
   assign soundFileAmplitudes [85] = 8'd133;
   assign soundFileAmplitudes [86] = 8'd139;
   assign soundFileAmplitudes [87] = 8'd141;
   assign soundFileAmplitudes [88] = 8'd149;
   assign soundFileAmplitudes [89] = 8'd115;
   assign soundFileAmplitudes [90] = 8'd118;
   assign soundFileAmplitudes [91] = 8'd131;
   assign soundFileAmplitudes [92] = 8'd120;
   assign soundFileAmplitudes [93] = 8'd125;
   assign soundFileAmplitudes [94] = 8'd121;
   assign soundFileAmplitudes [95] = 8'd115;
   assign soundFileAmplitudes [96] = 8'd114;
   assign soundFileAmplitudes [97] = 8'd112;
   assign soundFileAmplitudes [98] = 8'd102;
   assign soundFileAmplitudes [99] = 8'd108;
   assign soundFileAmplitudes [100] = 8'd127;
   assign soundFileAmplitudes [101] = 8'd133;
   assign soundFileAmplitudes [102] = 8'd131;
   assign soundFileAmplitudes [103] = 8'd115;
   assign soundFileAmplitudes [104] = 8'd114;
   assign soundFileAmplitudes [105] = 8'd130;
   assign soundFileAmplitudes [106] = 8'd128;
   assign soundFileAmplitudes [107] = 8'd143;
   assign soundFileAmplitudes [108] = 8'd139;
   assign soundFileAmplitudes [109] = 8'd147;
   assign soundFileAmplitudes [110] = 8'd137;
   assign soundFileAmplitudes [111] = 8'd111;
   assign soundFileAmplitudes [112] = 8'd125;
   assign soundFileAmplitudes [113] = 8'd142;
   assign soundFileAmplitudes [114] = 8'd151;
   assign soundFileAmplitudes [115] = 8'd142;
   assign soundFileAmplitudes [116] = 8'd138;
   assign soundFileAmplitudes [117] = 8'd137;
   assign soundFileAmplitudes [118] = 8'd131;
   assign soundFileAmplitudes [119] = 8'd114;
   assign soundFileAmplitudes [120] = 8'd121;
   assign soundFileAmplitudes [121] = 8'd133;
   assign soundFileAmplitudes [122] = 8'd136;
   assign soundFileAmplitudes [123] = 8'd126;
   assign soundFileAmplitudes [124] = 8'd123;
   assign soundFileAmplitudes [125] = 8'd120;
   assign soundFileAmplitudes [126] = 8'd120;
   assign soundFileAmplitudes [127] = 8'd133;
   assign soundFileAmplitudes [128] = 8'd132;
   assign soundFileAmplitudes [129] = 8'd126;
   assign soundFileAmplitudes [130] = 8'd117;
   assign soundFileAmplitudes [131] = 8'd110;
   assign soundFileAmplitudes [132] = 8'd101;
   assign soundFileAmplitudes [133] = 8'd107;
   assign soundFileAmplitudes [134] = 8'd113;
   assign soundFileAmplitudes [135] = 8'd125;
   assign soundFileAmplitudes [136] = 8'd123;
   assign soundFileAmplitudes [137] = 8'd123;
   assign soundFileAmplitudes [138] = 8'd122;
   assign soundFileAmplitudes [139] = 8'd130;
   assign soundFileAmplitudes [140] = 8'd144;
   assign soundFileAmplitudes [141] = 8'd141;
   assign soundFileAmplitudes [142] = 8'd143;
   assign soundFileAmplitudes [143] = 8'd142;
   assign soundFileAmplitudes [144] = 8'd146;
   assign soundFileAmplitudes [145] = 8'd130;
   assign soundFileAmplitudes [146] = 8'd122;
   assign soundFileAmplitudes [147] = 8'd138;
   assign soundFileAmplitudes [148] = 8'd145;
   assign soundFileAmplitudes [149] = 8'd135;
   assign soundFileAmplitudes [150] = 8'd116;
   assign soundFileAmplitudes [151] = 8'd117;
   assign soundFileAmplitudes [152] = 8'd124;
   assign soundFileAmplitudes [153] = 8'd127;
   assign soundFileAmplitudes [154] = 8'd121;
   assign soundFileAmplitudes [155] = 8'd116;
   assign soundFileAmplitudes [156] = 8'd129;
   assign soundFileAmplitudes [157] = 8'd136;
   assign soundFileAmplitudes [158] = 8'd148;
   assign soundFileAmplitudes [159] = 8'd131;
   assign soundFileAmplitudes [160] = 8'd114;
   assign soundFileAmplitudes [161] = 8'd119;
   assign soundFileAmplitudes [162] = 8'd122;
   assign soundFileAmplitudes [163] = 8'd129;
   assign soundFileAmplitudes [164] = 8'd113;
   assign soundFileAmplitudes [165] = 8'd102;
   assign soundFileAmplitudes [166] = 8'd94;
   assign soundFileAmplitudes [167] = 8'd87;
   assign soundFileAmplitudes [168] = 8'd103;
   assign soundFileAmplitudes [169] = 8'd128;
   assign soundFileAmplitudes [170] = 8'd144;
   assign soundFileAmplitudes [171] = 8'd149;
   assign soundFileAmplitudes [172] = 8'd139;
   assign soundFileAmplitudes [173] = 8'd132;
   assign soundFileAmplitudes [174] = 8'd145;
   assign soundFileAmplitudes [175] = 8'd149;
   assign soundFileAmplitudes [176] = 8'd140;
   assign soundFileAmplitudes [177] = 8'd134;
   assign soundFileAmplitudes [178] = 8'd129;
   assign soundFileAmplitudes [179] = 8'd129;
   assign soundFileAmplitudes [180] = 8'd105;
   assign soundFileAmplitudes [181] = 8'd104;
   assign soundFileAmplitudes [182] = 8'd124;
   assign soundFileAmplitudes [183] = 8'd125;
   assign soundFileAmplitudes [184] = 8'd121;
   assign soundFileAmplitudes [185] = 8'd107;
   assign soundFileAmplitudes [186] = 8'd114;
   assign soundFileAmplitudes [187] = 8'd141;
   assign soundFileAmplitudes [188] = 8'd147;
   assign soundFileAmplitudes [189] = 8'd141;
   assign soundFileAmplitudes [190] = 8'd130;
   assign soundFileAmplitudes [191] = 8'd120;
   assign soundFileAmplitudes [192] = 8'd132;
   assign soundFileAmplitudes [193] = 8'd133;
   assign soundFileAmplitudes [194] = 8'd128;
   assign soundFileAmplitudes [195] = 8'd122;
   assign soundFileAmplitudes [196] = 8'd121;
   assign soundFileAmplitudes [197] = 8'd115;
   assign soundFileAmplitudes [198] = 8'd103;
   assign soundFileAmplitudes [199] = 8'd118;
   assign soundFileAmplitudes [200] = 8'd123;
   assign soundFileAmplitudes [201] = 8'd123;
   assign soundFileAmplitudes [202] = 8'd117;
   assign soundFileAmplitudes [203] = 8'd116;
   assign soundFileAmplitudes [204] = 8'd131;
   assign soundFileAmplitudes [205] = 8'd153;
   assign soundFileAmplitudes [206] = 8'd152;
   assign soundFileAmplitudes [207] = 8'd139;
   assign soundFileAmplitudes [208] = 8'd134;
   assign soundFileAmplitudes [209] = 8'd141;
   assign soundFileAmplitudes [210] = 8'd145;
   assign soundFileAmplitudes [211] = 8'd121;
   assign soundFileAmplitudes [212] = 8'd116;
   assign soundFileAmplitudes [213] = 8'd116;
   assign soundFileAmplitudes [214] = 8'd109;
   assign soundFileAmplitudes [215] = 8'd94;
   assign soundFileAmplitudes [216] = 8'd94;
   assign soundFileAmplitudes [217] = 8'd117;
   assign soundFileAmplitudes [218] = 8'd124;
   assign soundFileAmplitudes [219] = 8'd131;
   assign soundFileAmplitudes [220] = 8'd135;
   assign soundFileAmplitudes [221] = 8'd138;
   assign soundFileAmplitudes [222] = 8'd139;
   assign soundFileAmplitudes [223] = 8'd144;
   assign soundFileAmplitudes [224] = 8'd141;
   assign soundFileAmplitudes [225] = 8'd135;
   assign soundFileAmplitudes [226] = 8'd140;
   assign soundFileAmplitudes [227] = 8'd129;
   assign soundFileAmplitudes [228] = 8'd115;
   assign soundFileAmplitudes [229] = 8'd112;
   assign soundFileAmplitudes [230] = 8'd121;
   assign soundFileAmplitudes [231] = 8'd129;
   assign soundFileAmplitudes [232] = 8'd129;
   assign soundFileAmplitudes [233] = 8'd127;
   assign soundFileAmplitudes [234] = 8'd124;
   assign soundFileAmplitudes [235] = 8'd123;
   assign soundFileAmplitudes [236] = 8'd130;
   assign soundFileAmplitudes [237] = 8'd123;
   assign soundFileAmplitudes [238] = 8'd126;
   assign soundFileAmplitudes [239] = 8'd142;
   assign soundFileAmplitudes [240] = 8'd145;
   assign soundFileAmplitudes [241] = 8'd138;
   assign soundFileAmplitudes [242] = 8'd113;
   assign soundFileAmplitudes [243] = 8'd118;
   assign soundFileAmplitudes [244] = 8'd134;
   assign soundFileAmplitudes [245] = 8'd140;
   assign soundFileAmplitudes [246] = 8'd133;
   assign soundFileAmplitudes [247] = 8'd118;
   assign soundFileAmplitudes [248] = 8'd116;
   assign soundFileAmplitudes [249] = 8'd125;
   assign soundFileAmplitudes [250] = 8'd126;
   assign soundFileAmplitudes [251] = 8'd122;
   assign soundFileAmplitudes [252] = 8'd113;
   assign soundFileAmplitudes [253] = 8'd110;
   assign soundFileAmplitudes [254] = 8'd127;
   assign soundFileAmplitudes [255] = 8'd136;
   assign soundFileAmplitudes [256] = 8'd127;
   assign soundFileAmplitudes [257] = 8'd125;
   assign soundFileAmplitudes [258] = 8'd117;
   assign soundFileAmplitudes [259] = 8'd105;
   assign soundFileAmplitudes [260] = 8'd119;
   assign soundFileAmplitudes [261] = 8'd132;
   assign soundFileAmplitudes [262] = 8'd139;
   assign soundFileAmplitudes [263] = 8'd147;
   assign soundFileAmplitudes [264] = 8'd138;
   assign soundFileAmplitudes [265] = 8'd130;
   assign soundFileAmplitudes [266] = 8'd133;
   assign soundFileAmplitudes [267] = 8'd150;
   assign soundFileAmplitudes [268] = 8'd143;
   assign soundFileAmplitudes [269] = 8'd136;
   assign soundFileAmplitudes [270] = 8'd132;
   assign soundFileAmplitudes [271] = 8'd129;
   assign soundFileAmplitudes [272] = 8'd130;
   assign soundFileAmplitudes [273] = 8'd97;
   assign soundFileAmplitudes [274] = 8'd105;
   assign soundFileAmplitudes [275] = 8'd122;
   assign soundFileAmplitudes [276] = 8'd123;
   assign soundFileAmplitudes [277] = 8'd123;
   assign soundFileAmplitudes [278] = 8'd112;
   assign soundFileAmplitudes [279] = 8'd125;
   assign soundFileAmplitudes [280] = 8'd140;
   assign soundFileAmplitudes [281] = 8'd149;
   assign soundFileAmplitudes [282] = 8'd146;
   assign soundFileAmplitudes [283] = 8'd132;
   assign soundFileAmplitudes [284] = 8'd134;
   assign soundFileAmplitudes [285] = 8'd124;
   assign soundFileAmplitudes [286] = 8'd109;
   assign soundFileAmplitudes [287] = 8'd114;
   assign soundFileAmplitudes [288] = 8'd115;
   assign soundFileAmplitudes [289] = 8'd117;
   assign soundFileAmplitudes [290] = 8'd100;
   assign soundFileAmplitudes [291] = 8'd100;
   assign soundFileAmplitudes [292] = 8'd115;
   assign soundFileAmplitudes [293] = 8'd122;
   assign soundFileAmplitudes [294] = 8'd132;
   assign soundFileAmplitudes [295] = 8'd124;
   assign soundFileAmplitudes [296] = 8'd127;
   assign soundFileAmplitudes [297] = 8'd137;
   assign soundFileAmplitudes [298] = 8'd153;
   assign soundFileAmplitudes [299] = 8'd154;
   assign soundFileAmplitudes [300] = 8'd146;
   assign soundFileAmplitudes [301] = 8'd143;
   assign soundFileAmplitudes [302] = 8'd146;
   assign soundFileAmplitudes [303] = 8'd150;
   assign soundFileAmplitudes [304] = 8'd121;
   assign soundFileAmplitudes [305] = 8'd105;
   assign soundFileAmplitudes [306] = 8'd107;
   assign soundFileAmplitudes [307] = 8'd108;
   assign soundFileAmplitudes [308] = 8'd112;
   assign soundFileAmplitudes [309] = 8'd116;
   assign soundFileAmplitudes [310] = 8'd120;
   assign soundFileAmplitudes [311] = 8'd128;
   assign soundFileAmplitudes [312] = 8'd134;
   assign soundFileAmplitudes [313] = 8'd129;
   assign soundFileAmplitudes [314] = 8'd129;
   assign soundFileAmplitudes [315] = 8'd144;
   assign soundFileAmplitudes [316] = 8'd145;
   assign soundFileAmplitudes [317] = 8'd142;
   assign soundFileAmplitudes [318] = 8'd138;
   assign soundFileAmplitudes [319] = 8'd126;
   assign soundFileAmplitudes [320] = 8'd113;
   assign soundFileAmplitudes [321] = 8'd90;
   assign soundFileAmplitudes [322] = 8'd98;
   assign soundFileAmplitudes [323] = 8'd118;
   assign soundFileAmplitudes [324] = 8'd122;
   assign soundFileAmplitudes [325] = 8'd120;
   assign soundFileAmplitudes [326] = 8'd111;
   assign soundFileAmplitudes [327] = 8'd110;
   assign soundFileAmplitudes [328] = 8'd113;
   assign soundFileAmplitudes [329] = 8'd113;
   assign soundFileAmplitudes [330] = 8'd124;
   assign soundFileAmplitudes [331] = 8'd136;
   assign soundFileAmplitudes [332] = 8'd142;
   assign soundFileAmplitudes [333] = 8'd147;
   assign soundFileAmplitudes [334] = 8'd138;
   assign soundFileAmplitudes [335] = 8'd126;
   assign soundFileAmplitudes [336] = 8'd121;
   assign soundFileAmplitudes [337] = 8'd135;
   assign soundFileAmplitudes [338] = 8'd142;
   assign soundFileAmplitudes [339] = 8'd135;
   assign soundFileAmplitudes [340] = 8'd125;
   assign soundFileAmplitudes [341] = 8'd120;
   assign soundFileAmplitudes [342] = 8'd127;
   assign soundFileAmplitudes [343] = 8'd134;
   assign soundFileAmplitudes [344] = 8'd134;
   assign soundFileAmplitudes [345] = 8'd131;
   assign soundFileAmplitudes [346] = 8'd136;
   assign soundFileAmplitudes [347] = 8'd132;
   assign soundFileAmplitudes [348] = 8'd124;
   assign soundFileAmplitudes [349] = 8'd128;
   assign soundFileAmplitudes [350] = 8'd132;
   assign soundFileAmplitudes [351] = 8'd133;
   assign soundFileAmplitudes [352] = 8'd127;
   assign soundFileAmplitudes [353] = 8'd123;
   assign soundFileAmplitudes [354] = 8'd127;
   assign soundFileAmplitudes [355] = 8'd116;
   assign soundFileAmplitudes [356] = 8'd115;
   assign soundFileAmplitudes [357] = 8'd126;
   assign soundFileAmplitudes [358] = 8'd123;
   assign soundFileAmplitudes [359] = 8'd116;
   assign soundFileAmplitudes [360] = 8'd120;
   assign soundFileAmplitudes [361] = 8'd111;
   assign soundFileAmplitudes [362] = 8'd124;
   assign soundFileAmplitudes [363] = 8'd123;
   assign soundFileAmplitudes [364] = 8'd105;
   assign soundFileAmplitudes [365] = 8'd105;
   assign soundFileAmplitudes [366] = 8'd105;
   assign soundFileAmplitudes [367] = 8'd120;
   assign soundFileAmplitudes [368] = 8'd135;
   assign soundFileAmplitudes [369] = 8'd140;
   assign soundFileAmplitudes [370] = 8'd130;
   assign soundFileAmplitudes [371] = 8'd135;
   assign soundFileAmplitudes [372] = 8'd141;
   assign soundFileAmplitudes [373] = 8'd146;
   assign soundFileAmplitudes [374] = 8'd154;
   assign soundFileAmplitudes [375] = 8'd145;
   assign soundFileAmplitudes [376] = 8'd127;
   assign soundFileAmplitudes [377] = 8'd127;
   assign soundFileAmplitudes [378] = 8'd133;
   assign soundFileAmplitudes [379] = 8'd133;
   assign soundFileAmplitudes [380] = 8'd132;
   assign soundFileAmplitudes [381] = 8'd126;
   assign soundFileAmplitudes [382] = 8'd123;
   assign soundFileAmplitudes [383] = 8'd111;
   assign soundFileAmplitudes [384] = 8'd115;
   assign soundFileAmplitudes [385] = 8'd130;
   assign soundFileAmplitudes [386] = 8'd141;
   assign soundFileAmplitudes [387] = 8'd150;
   assign soundFileAmplitudes [388] = 8'd139;
   assign soundFileAmplitudes [389] = 8'd131;
   assign soundFileAmplitudes [390] = 8'd123;
   assign soundFileAmplitudes [391] = 8'd120;
   assign soundFileAmplitudes [392] = 8'd128;
   assign soundFileAmplitudes [393] = 8'd134;
   assign soundFileAmplitudes [394] = 8'd125;
   assign soundFileAmplitudes [395] = 8'd112;
   assign soundFileAmplitudes [396] = 8'd95;
   assign soundFileAmplitudes [397] = 8'd96;
   assign soundFileAmplitudes [398] = 8'd99;
   assign soundFileAmplitudes [399] = 8'd100;
   assign soundFileAmplitudes [400] = 8'd113;
   assign soundFileAmplitudes [401] = 8'd112;
   assign soundFileAmplitudes [402] = 8'd127;
   assign soundFileAmplitudes [403] = 8'd133;
   assign soundFileAmplitudes [404] = 8'd134;
   assign soundFileAmplitudes [405] = 8'd149;
   assign soundFileAmplitudes [406] = 8'd149;
   assign soundFileAmplitudes [407] = 8'd143;
   assign soundFileAmplitudes [408] = 8'd154;
   assign soundFileAmplitudes [409] = 8'd155;
   assign soundFileAmplitudes [410] = 8'd143;
   assign soundFileAmplitudes [411] = 8'd128;
   assign soundFileAmplitudes [412] = 8'd122;
   assign soundFileAmplitudes [413] = 8'd119;
   assign soundFileAmplitudes [414] = 8'd116;
   assign soundFileAmplitudes [415] = 8'd132;
   assign soundFileAmplitudes [416] = 8'd146;
   assign soundFileAmplitudes [417] = 8'd140;
   assign soundFileAmplitudes [418] = 8'd130;
   assign soundFileAmplitudes [419] = 8'd120;
   assign soundFileAmplitudes [420] = 8'd130;
   assign soundFileAmplitudes [421] = 8'd149;
   assign soundFileAmplitudes [422] = 8'd146;
   assign soundFileAmplitudes [423] = 8'd144;
   assign soundFileAmplitudes [424] = 8'd132;
   assign soundFileAmplitudes [425] = 8'd111;
   assign soundFileAmplitudes [426] = 8'd86;
   assign soundFileAmplitudes [427] = 8'd94;
   assign soundFileAmplitudes [428] = 8'd104;
   assign soundFileAmplitudes [429] = 8'd106;
   assign soundFileAmplitudes [430] = 8'd104;
   assign soundFileAmplitudes [431] = 8'd100;
   assign soundFileAmplitudes [432] = 8'd107;
   assign soundFileAmplitudes [433] = 8'd108;
   assign soundFileAmplitudes [434] = 8'd125;
   assign soundFileAmplitudes [435] = 8'd134;
   assign soundFileAmplitudes [436] = 8'd126;
   assign soundFileAmplitudes [437] = 8'd135;
   assign soundFileAmplitudes [438] = 8'd147;
   assign soundFileAmplitudes [439] = 8'd143;
   assign soundFileAmplitudes [440] = 8'd136;
   assign soundFileAmplitudes [441] = 8'd128;
   assign soundFileAmplitudes [442] = 8'd130;
   assign soundFileAmplitudes [443] = 8'd128;
   assign soundFileAmplitudes [444] = 8'd125;
   assign soundFileAmplitudes [445] = 8'd133;
   assign soundFileAmplitudes [446] = 8'd138;
   assign soundFileAmplitudes [447] = 8'd133;
   assign soundFileAmplitudes [448] = 8'd138;
   assign soundFileAmplitudes [449] = 8'd142;
   assign soundFileAmplitudes [450] = 8'd155;
   assign soundFileAmplitudes [451] = 8'd152;
   assign soundFileAmplitudes [452] = 8'd141;
   assign soundFileAmplitudes [453] = 8'd142;
   assign soundFileAmplitudes [454] = 8'd138;
   assign soundFileAmplitudes [455] = 8'd128;
   assign soundFileAmplitudes [456] = 8'd107;
   assign soundFileAmplitudes [457] = 8'd113;
   assign soundFileAmplitudes [458] = 8'd112;
   assign soundFileAmplitudes [459] = 8'd105;
   assign soundFileAmplitudes [460] = 8'd101;
   assign soundFileAmplitudes [461] = 8'd87;
   assign soundFileAmplitudes [462] = 8'd90;
   assign soundFileAmplitudes [463] = 8'd109;
   assign soundFileAmplitudes [464] = 8'd116;
   assign soundFileAmplitudes [465] = 8'd117;
   assign soundFileAmplitudes [466] = 8'd116;
   assign soundFileAmplitudes [467] = 8'd125;
   assign soundFileAmplitudes [468] = 8'd138;
   assign soundFileAmplitudes [469] = 8'd136;
   assign soundFileAmplitudes [470] = 8'd131;
   assign soundFileAmplitudes [471] = 8'd129;
   assign soundFileAmplitudes [472] = 8'd128;
   assign soundFileAmplitudes [473] = 8'd126;
   assign soundFileAmplitudes [474] = 8'd122;
   assign soundFileAmplitudes [475] = 8'd127;
   assign soundFileAmplitudes [476] = 8'd142;
   assign soundFileAmplitudes [477] = 8'd147;
   assign soundFileAmplitudes [478] = 8'd152;
   assign soundFileAmplitudes [479] = 8'd150;
   assign soundFileAmplitudes [480] = 8'd153;
   assign soundFileAmplitudes [481] = 8'd147;
   assign soundFileAmplitudes [482] = 8'd133;
   assign soundFileAmplitudes [483] = 8'd134;
   assign soundFileAmplitudes [484] = 8'd137;
   assign soundFileAmplitudes [485] = 8'd129;
   assign soundFileAmplitudes [486] = 8'd107;
   assign soundFileAmplitudes [487] = 8'd111;
   assign soundFileAmplitudes [488] = 8'd118;
   assign soundFileAmplitudes [489] = 8'd108;
   assign soundFileAmplitudes [490] = 8'd108;
   assign soundFileAmplitudes [491] = 8'd111;
   assign soundFileAmplitudes [492] = 8'd113;
   assign soundFileAmplitudes [493] = 8'd122;
   assign soundFileAmplitudes [494] = 8'd133;
   assign soundFileAmplitudes [495] = 8'd134;
   assign soundFileAmplitudes [496] = 8'd118;
   assign soundFileAmplitudes [497] = 8'd116;
   assign soundFileAmplitudes [498] = 8'd121;
   assign soundFileAmplitudes [499] = 8'd119;
   assign soundFileAmplitudes [500] = 8'd121;
   assign soundFileAmplitudes [501] = 8'd121;
   assign soundFileAmplitudes [502] = 8'd119;
   assign soundFileAmplitudes [503] = 8'd107;
   assign soundFileAmplitudes [504] = 8'd99;
   assign soundFileAmplitudes [505] = 8'd112;
   assign soundFileAmplitudes [506] = 8'd128;
   assign soundFileAmplitudes [507] = 8'd138;
   assign soundFileAmplitudes [508] = 8'd141;
   assign soundFileAmplitudes [509] = 8'd143;
   assign soundFileAmplitudes [510] = 8'd153;
   assign soundFileAmplitudes [511] = 8'd167;
   assign soundFileAmplitudes [512] = 8'd159;
   assign soundFileAmplitudes [513] = 8'd155;
   assign soundFileAmplitudes [514] = 8'd154;
   assign soundFileAmplitudes [515] = 8'd152;
   assign soundFileAmplitudes [516] = 8'd133;
   assign soundFileAmplitudes [517] = 8'd103;
   assign soundFileAmplitudes [518] = 8'd107;
   assign soundFileAmplitudes [519] = 8'd120;
   assign soundFileAmplitudes [520] = 8'd114;
   assign soundFileAmplitudes [521] = 8'd102;
   assign soundFileAmplitudes [522] = 8'd101;
   assign soundFileAmplitudes [523] = 8'd110;
   assign soundFileAmplitudes [524] = 8'd122;
   assign soundFileAmplitudes [525] = 8'd133;
   assign soundFileAmplitudes [526] = 8'd142;
   assign soundFileAmplitudes [527] = 8'd140;
   assign soundFileAmplitudes [528] = 8'd138;
   assign soundFileAmplitudes [529] = 8'd136;
   assign soundFileAmplitudes [530] = 8'd141;
   assign soundFileAmplitudes [531] = 8'd134;
   assign soundFileAmplitudes [532] = 8'd114;
   assign soundFileAmplitudes [533] = 8'd114;
   assign soundFileAmplitudes [534] = 8'd104;
   assign soundFileAmplitudes [535] = 8'd103;
   assign soundFileAmplitudes [536] = 8'd121;
   assign soundFileAmplitudes [537] = 8'd116;
   assign soundFileAmplitudes [538] = 8'd111;
   assign soundFileAmplitudes [539] = 8'd110;
   assign soundFileAmplitudes [540] = 8'd119;
   assign soundFileAmplitudes [541] = 8'd137;
   assign soundFileAmplitudes [542] = 8'd148;
   assign soundFileAmplitudes [543] = 8'd151;
   assign soundFileAmplitudes [544] = 8'd146;
   assign soundFileAmplitudes [545] = 8'd148;
   assign soundFileAmplitudes [546] = 8'd156;
   assign soundFileAmplitudes [547] = 8'd144;
   assign soundFileAmplitudes [548] = 8'd121;
   assign soundFileAmplitudes [549] = 8'd128;
   assign soundFileAmplitudes [550] = 8'd139;
   assign soundFileAmplitudes [551] = 8'd132;
   assign soundFileAmplitudes [552] = 8'd113;
   assign soundFileAmplitudes [553] = 8'd104;
   assign soundFileAmplitudes [554] = 8'd114;
   assign soundFileAmplitudes [555] = 8'd125;
   assign soundFileAmplitudes [556] = 8'd130;
   assign soundFileAmplitudes [557] = 8'd125;
   assign soundFileAmplitudes [558] = 8'd123;
   assign soundFileAmplitudes [559] = 8'd122;
   assign soundFileAmplitudes [560] = 8'd122;
   assign soundFileAmplitudes [561] = 8'd128;
   assign soundFileAmplitudes [562] = 8'd125;
   assign soundFileAmplitudes [563] = 8'd124;
   assign soundFileAmplitudes [564] = 8'd118;
   assign soundFileAmplitudes [565] = 8'd110;
   assign soundFileAmplitudes [566] = 8'd113;
   assign soundFileAmplitudes [567] = 8'd119;
   assign soundFileAmplitudes [568] = 8'd132;
   assign soundFileAmplitudes [569] = 8'd117;
   assign soundFileAmplitudes [570] = 8'd111;
   assign soundFileAmplitudes [571] = 8'd121;
   assign soundFileAmplitudes [572] = 8'd128;
   assign soundFileAmplitudes [573] = 8'd143;
   assign soundFileAmplitudes [574] = 8'd123;
   assign soundFileAmplitudes [575] = 8'd111;
   assign soundFileAmplitudes [576] = 8'd135;
   assign soundFileAmplitudes [577] = 8'd146;
   assign soundFileAmplitudes [578] = 8'd142;
   assign soundFileAmplitudes [579] = 8'd117;
   assign soundFileAmplitudes [580] = 8'd114;
   assign soundFileAmplitudes [581] = 8'd138;
   assign soundFileAmplitudes [582] = 8'd135;
   assign soundFileAmplitudes [583] = 8'd131;
   assign soundFileAmplitudes [584] = 8'd135;
   assign soundFileAmplitudes [585] = 8'd142;
   assign soundFileAmplitudes [586] = 8'd138;
   assign soundFileAmplitudes [587] = 8'd121;
   assign soundFileAmplitudes [588] = 8'd113;
   assign soundFileAmplitudes [589] = 8'd120;
   assign soundFileAmplitudes [590] = 8'd135;
   assign soundFileAmplitudes [591] = 8'd139;
   assign soundFileAmplitudes [592] = 8'd131;
   assign soundFileAmplitudes [593] = 8'd122;
   assign soundFileAmplitudes [594] = 8'd122;
   assign soundFileAmplitudes [595] = 8'd114;
   assign soundFileAmplitudes [596] = 8'd122;
   assign soundFileAmplitudes [597] = 8'd130;
   assign soundFileAmplitudes [598] = 8'd135;
   assign soundFileAmplitudes [599] = 8'd138;
   assign soundFileAmplitudes [600] = 8'd133;
   assign soundFileAmplitudes [601] = 8'd118;
   assign soundFileAmplitudes [602] = 8'd105;
   assign soundFileAmplitudes [603] = 8'd113;
   assign soundFileAmplitudes [604] = 8'd112;
   assign soundFileAmplitudes [605] = 8'd112;
   assign soundFileAmplitudes [606] = 8'd99;
   assign soundFileAmplitudes [607] = 8'd114;
   assign soundFileAmplitudes [608] = 8'd135;
   assign soundFileAmplitudes [609] = 8'd134;
   assign soundFileAmplitudes [610] = 8'd109;
   assign soundFileAmplitudes [611] = 8'd100;
   assign soundFileAmplitudes [612] = 8'd131;
   assign soundFileAmplitudes [613] = 8'd141;
   assign soundFileAmplitudes [614] = 8'd142;
   assign soundFileAmplitudes [615] = 8'd144;
   assign soundFileAmplitudes [616] = 8'd155;
   assign soundFileAmplitudes [617] = 8'd156;
   assign soundFileAmplitudes [618] = 8'd150;
   assign soundFileAmplitudes [619] = 8'd142;
   assign soundFileAmplitudes [620] = 8'd136;
   assign soundFileAmplitudes [621] = 8'd119;
   assign soundFileAmplitudes [622] = 8'd103;
   assign soundFileAmplitudes [623] = 8'd107;
   assign soundFileAmplitudes [624] = 8'd111;
   assign soundFileAmplitudes [625] = 8'd106;
   assign soundFileAmplitudes [626] = 8'd106;
   assign soundFileAmplitudes [627] = 8'd126;
   assign soundFileAmplitudes [628] = 8'd138;
   assign soundFileAmplitudes [629] = 8'd142;
   assign soundFileAmplitudes [630] = 8'd142;
   assign soundFileAmplitudes [631] = 8'd146;
   assign soundFileAmplitudes [632] = 8'd142;
   assign soundFileAmplitudes [633] = 8'd138;
   assign soundFileAmplitudes [634] = 8'd133;
   assign soundFileAmplitudes [635] = 8'd136;
   assign soundFileAmplitudes [636] = 8'd115;
   assign soundFileAmplitudes [637] = 8'd91;
   assign soundFileAmplitudes [638] = 8'd99;
   assign soundFileAmplitudes [639] = 8'd100;
   assign soundFileAmplitudes [640] = 8'd97;
   assign soundFileAmplitudes [641] = 8'd81;
   assign soundFileAmplitudes [642] = 8'd98;
   assign soundFileAmplitudes [643] = 8'd120;
   assign soundFileAmplitudes [644] = 8'd126;
   assign soundFileAmplitudes [645] = 8'd131;
   assign soundFileAmplitudes [646] = 8'd139;
   assign soundFileAmplitudes [647] = 8'd161;
   assign soundFileAmplitudes [648] = 8'd175;
   assign soundFileAmplitudes [649] = 8'd172;
   assign soundFileAmplitudes [650] = 8'd171;
   assign soundFileAmplitudes [651] = 8'd158;
   assign soundFileAmplitudes [652] = 8'd142;
   assign soundFileAmplitudes [653] = 8'd137;
   assign soundFileAmplitudes [654] = 8'd125;
   assign soundFileAmplitudes [655] = 8'd115;
   assign soundFileAmplitudes [656] = 8'd94;
   assign soundFileAmplitudes [657] = 8'd92;
   assign soundFileAmplitudes [658] = 8'd108;
   assign soundFileAmplitudes [659] = 8'd120;
   assign soundFileAmplitudes [660] = 8'd131;
   assign soundFileAmplitudes [661] = 8'd132;
   assign soundFileAmplitudes [662] = 8'd132;
   assign soundFileAmplitudes [663] = 8'd136;
   assign soundFileAmplitudes [664] = 8'd136;
   assign soundFileAmplitudes [665] = 8'd142;
   assign soundFileAmplitudes [666] = 8'd146;
   assign soundFileAmplitudes [667] = 8'd129;
   assign soundFileAmplitudes [668] = 8'd131;
   assign soundFileAmplitudes [669] = 8'd136;
   assign soundFileAmplitudes [670] = 8'd135;
   assign soundFileAmplitudes [671] = 8'd104;
   assign soundFileAmplitudes [672] = 8'd67;
   assign soundFileAmplitudes [673] = 8'd75;
   assign soundFileAmplitudes [674] = 8'd87;
   assign soundFileAmplitudes [675] = 8'd103;
   assign soundFileAmplitudes [676] = 8'd117;
   assign soundFileAmplitudes [677] = 8'd125;
   assign soundFileAmplitudes [678] = 8'd130;
   assign soundFileAmplitudes [679] = 8'd137;
   assign soundFileAmplitudes [680] = 8'd140;
   assign soundFileAmplitudes [681] = 8'd155;
   assign soundFileAmplitudes [682] = 8'd167;
   assign soundFileAmplitudes [683] = 8'd163;
   assign soundFileAmplitudes [684] = 8'd148;
   assign soundFileAmplitudes [685] = 8'd141;
   assign soundFileAmplitudes [686] = 8'd133;
   assign soundFileAmplitudes [687] = 8'd123;
   assign soundFileAmplitudes [688] = 8'd137;
   assign soundFileAmplitudes [689] = 8'd133;
   assign soundFileAmplitudes [690] = 8'd123;
   assign soundFileAmplitudes [691] = 8'd116;
   assign soundFileAmplitudes [692] = 8'd109;
   assign soundFileAmplitudes [693] = 8'd114;
   assign soundFileAmplitudes [694] = 8'd122;
   assign soundFileAmplitudes [695] = 8'd132;
   assign soundFileAmplitudes [696] = 8'd131;
   assign soundFileAmplitudes [697] = 8'd117;
   assign soundFileAmplitudes [698] = 8'd108;
   assign soundFileAmplitudes [699] = 8'd114;
   assign soundFileAmplitudes [700] = 8'd130;
   assign soundFileAmplitudes [701] = 8'd127;
   assign soundFileAmplitudes [702] = 8'd105;
   assign soundFileAmplitudes [703] = 8'd115;
   assign soundFileAmplitudes [704] = 8'd133;
   assign soundFileAmplitudes [705] = 8'd129;
   assign soundFileAmplitudes [706] = 8'd113;
   assign soundFileAmplitudes [707] = 8'd115;
   assign soundFileAmplitudes [708] = 8'd128;
   assign soundFileAmplitudes [709] = 8'd127;
   assign soundFileAmplitudes [710] = 8'd130;
   assign soundFileAmplitudes [711] = 8'd128;
   assign soundFileAmplitudes [712] = 8'd134;
   assign soundFileAmplitudes [713] = 8'd137;
   assign soundFileAmplitudes [714] = 8'd131;
   assign soundFileAmplitudes [715] = 8'd138;
   assign soundFileAmplitudes [716] = 8'd137;
   assign soundFileAmplitudes [717] = 8'd132;
   assign soundFileAmplitudes [718] = 8'd134;
   assign soundFileAmplitudes [719] = 8'd134;
   assign soundFileAmplitudes [720] = 8'd138;
   assign soundFileAmplitudes [721] = 8'd133;
   assign soundFileAmplitudes [722] = 8'd131;
   assign soundFileAmplitudes [723] = 8'd135;
   assign soundFileAmplitudes [724] = 8'd129;
   assign soundFileAmplitudes [725] = 8'd122;
   assign soundFileAmplitudes [726] = 8'd124;
   assign soundFileAmplitudes [727] = 8'd119;
   assign soundFileAmplitudes [728] = 8'd115;
   assign soundFileAmplitudes [729] = 8'd109;
   assign soundFileAmplitudes [730] = 8'd104;
   assign soundFileAmplitudes [731] = 8'd121;
   assign soundFileAmplitudes [732] = 8'd116;
   assign soundFileAmplitudes [733] = 8'd101;
   assign soundFileAmplitudes [734] = 8'd94;
   assign soundFileAmplitudes [735] = 8'd110;
   assign soundFileAmplitudes [736] = 8'd126;
   assign soundFileAmplitudes [737] = 8'd125;
   assign soundFileAmplitudes [738] = 8'd124;
   assign soundFileAmplitudes [739] = 8'd127;
   assign soundFileAmplitudes [740] = 8'd147;
   assign soundFileAmplitudes [741] = 8'd153;
   assign soundFileAmplitudes [742] = 8'd140;
   assign soundFileAmplitudes [743] = 8'd128;
   assign soundFileAmplitudes [744] = 8'd132;
   assign soundFileAmplitudes [745] = 8'd138;
   assign soundFileAmplitudes [746] = 8'd134;
   assign soundFileAmplitudes [747] = 8'd126;
   assign soundFileAmplitudes [748] = 8'd112;
   assign soundFileAmplitudes [749] = 8'd112;
   assign soundFileAmplitudes [750] = 8'd133;
   assign soundFileAmplitudes [751] = 8'd149;
   assign soundFileAmplitudes [752] = 8'd151;
   assign soundFileAmplitudes [753] = 8'd139;
   assign soundFileAmplitudes [754] = 8'd127;
   assign soundFileAmplitudes [755] = 8'd130;
   assign soundFileAmplitudes [756] = 8'd134;
   assign soundFileAmplitudes [757] = 8'd138;
   assign soundFileAmplitudes [758] = 8'd142;
   assign soundFileAmplitudes [759] = 8'd130;
   assign soundFileAmplitudes [760] = 8'd113;
   assign soundFileAmplitudes [761] = 8'd109;
   assign soundFileAmplitudes [762] = 8'd122;
   assign soundFileAmplitudes [763] = 8'd122;
   assign soundFileAmplitudes [764] = 8'd107;
   assign soundFileAmplitudes [765] = 8'd100;
   assign soundFileAmplitudes [766] = 8'd110;
   assign soundFileAmplitudes [767] = 8'd115;
   assign soundFileAmplitudes [768] = 8'd116;
   assign soundFileAmplitudes [769] = 8'd132;
   assign soundFileAmplitudes [770] = 8'd142;
   assign soundFileAmplitudes [771] = 8'd144;
   assign soundFileAmplitudes [772] = 8'd137;
   assign soundFileAmplitudes [773] = 8'd133;
   assign soundFileAmplitudes [774] = 8'd136;
   assign soundFileAmplitudes [775] = 8'd132;
   assign soundFileAmplitudes [776] = 8'd121;
   assign soundFileAmplitudes [777] = 8'd113;
   assign soundFileAmplitudes [778] = 8'd107;
   assign soundFileAmplitudes [779] = 8'd100;
   assign soundFileAmplitudes [780] = 8'd107;
   assign soundFileAmplitudes [781] = 8'd116;
   assign soundFileAmplitudes [782] = 8'd124;
   assign soundFileAmplitudes [783] = 8'd127;
   assign soundFileAmplitudes [784] = 8'd131;
   assign soundFileAmplitudes [785] = 8'd133;
   assign soundFileAmplitudes [786] = 8'd141;
   assign soundFileAmplitudes [787] = 8'd149;
   assign soundFileAmplitudes [788] = 8'd154;
   assign soundFileAmplitudes [789] = 8'd142;
   assign soundFileAmplitudes [790] = 8'd136;
   assign soundFileAmplitudes [791] = 8'd144;
   assign soundFileAmplitudes [792] = 8'd143;
   assign soundFileAmplitudes [793] = 8'd134;
   assign soundFileAmplitudes [794] = 8'd107;
   assign soundFileAmplitudes [795] = 8'd96;
   assign soundFileAmplitudes [796] = 8'd109;
   assign soundFileAmplitudes [797] = 8'd116;
   assign soundFileAmplitudes [798] = 8'd117;
   assign soundFileAmplitudes [799] = 8'd128;
   assign soundFileAmplitudes [800] = 8'd145;
   assign soundFileAmplitudes [801] = 8'd149;
   assign soundFileAmplitudes [802] = 8'd141;
   assign soundFileAmplitudes [803] = 8'd137;
   assign soundFileAmplitudes [804] = 8'd130;
   assign soundFileAmplitudes [805] = 8'd141;
   assign soundFileAmplitudes [806] = 8'd136;
   assign soundFileAmplitudes [807] = 8'd124;
   assign soundFileAmplitudes [808] = 8'd116;
   assign soundFileAmplitudes [809] = 8'd110;
   assign soundFileAmplitudes [810] = 8'd114;
   assign soundFileAmplitudes [811] = 8'd103;
   assign soundFileAmplitudes [812] = 8'd108;
   assign soundFileAmplitudes [813] = 8'd106;
   assign soundFileAmplitudes [814] = 8'd107;
   assign soundFileAmplitudes [815] = 8'd125;
   assign soundFileAmplitudes [816] = 8'd131;
   assign soundFileAmplitudes [817] = 8'd138;
   assign soundFileAmplitudes [818] = 8'd135;
   assign soundFileAmplitudes [819] = 8'd124;
   assign soundFileAmplitudes [820] = 8'd137;
   assign soundFileAmplitudes [821] = 8'd141;
   assign soundFileAmplitudes [822] = 8'd142;
   assign soundFileAmplitudes [823] = 8'd131;
   assign soundFileAmplitudes [824] = 8'd114;
   assign soundFileAmplitudes [825] = 8'd129;
   assign soundFileAmplitudes [826] = 8'd132;
   assign soundFileAmplitudes [827] = 8'd129;
   assign soundFileAmplitudes [828] = 8'd126;
   assign soundFileAmplitudes [829] = 8'd125;
   assign soundFileAmplitudes [830] = 8'd127;
   assign soundFileAmplitudes [831] = 8'd129;
   assign soundFileAmplitudes [832] = 8'd126;
   assign soundFileAmplitudes [833] = 8'd127;
   assign soundFileAmplitudes [834] = 8'd137;
   assign soundFileAmplitudes [835] = 8'd142;
   assign soundFileAmplitudes [836] = 8'd136;
   assign soundFileAmplitudes [837] = 8'd123;
   assign soundFileAmplitudes [838] = 8'd114;
   assign soundFileAmplitudes [839] = 8'd116;
   assign soundFileAmplitudes [840] = 8'd115;
   assign soundFileAmplitudes [841] = 8'd121;
   assign soundFileAmplitudes [842] = 8'd130;
   assign soundFileAmplitudes [843] = 8'd131;
   assign soundFileAmplitudes [844] = 8'd126;
   assign soundFileAmplitudes [845] = 8'd101;
   assign soundFileAmplitudes [846] = 8'd102;
   assign soundFileAmplitudes [847] = 8'd109;
   assign soundFileAmplitudes [848] = 8'd118;
   assign soundFileAmplitudes [849] = 8'd130;
   assign soundFileAmplitudes [850] = 8'd118;
   assign soundFileAmplitudes [851] = 8'd121;
   assign soundFileAmplitudes [852] = 8'd126;
   assign soundFileAmplitudes [853] = 8'd128;
   assign soundFileAmplitudes [854] = 8'd126;
   assign soundFileAmplitudes [855] = 8'd113;
   assign soundFileAmplitudes [856] = 8'd127;
   assign soundFileAmplitudes [857] = 8'd148;
   assign soundFileAmplitudes [858] = 8'd147;
   assign soundFileAmplitudes [859] = 8'd138;
   assign soundFileAmplitudes [860] = 8'd138;
   assign soundFileAmplitudes [861] = 8'd145;
   assign soundFileAmplitudes [862] = 8'd149;
   assign soundFileAmplitudes [863] = 8'd145;
   assign soundFileAmplitudes [864] = 8'd133;
   assign soundFileAmplitudes [865] = 8'd124;
   assign soundFileAmplitudes [866] = 8'd115;
   assign soundFileAmplitudes [867] = 8'd113;
   assign soundFileAmplitudes [868] = 8'd117;
   assign soundFileAmplitudes [869] = 8'd124;
   assign soundFileAmplitudes [870] = 8'd113;
   assign soundFileAmplitudes [871] = 8'd103;
   assign soundFileAmplitudes [872] = 8'd112;
   assign soundFileAmplitudes [873] = 8'd128;
   assign soundFileAmplitudes [874] = 8'd147;
   assign soundFileAmplitudes [875] = 8'd146;
   assign soundFileAmplitudes [876] = 8'd144;
   assign soundFileAmplitudes [877] = 8'd139;
   assign soundFileAmplitudes [878] = 8'd132;
   assign soundFileAmplitudes [879] = 8'd126;
   assign soundFileAmplitudes [880] = 8'd117;
   assign soundFileAmplitudes [881] = 8'd112;
   assign soundFileAmplitudes [882] = 8'd109;
   assign soundFileAmplitudes [883] = 8'd103;
   assign soundFileAmplitudes [884] = 8'd107;
   assign soundFileAmplitudes [885] = 8'd114;
   assign soundFileAmplitudes [886] = 8'd101;
   assign soundFileAmplitudes [887] = 8'd96;
   assign soundFileAmplitudes [888] = 8'd105;
   assign soundFileAmplitudes [889] = 8'd121;
   assign soundFileAmplitudes [890] = 8'd138;
   assign soundFileAmplitudes [891] = 8'd150;
   assign soundFileAmplitudes [892] = 8'd153;
   assign soundFileAmplitudes [893] = 8'd149;
   assign soundFileAmplitudes [894] = 8'd144;
   assign soundFileAmplitudes [895] = 8'd145;
   assign soundFileAmplitudes [896] = 8'd150;
   assign soundFileAmplitudes [897] = 8'd151;
   assign soundFileAmplitudes [898] = 8'd142;
   assign soundFileAmplitudes [899] = 8'd125;
   assign soundFileAmplitudes [900] = 8'd109;
   assign soundFileAmplitudes [901] = 8'd107;
   assign soundFileAmplitudes [902] = 8'd109;
   assign soundFileAmplitudes [903] = 8'd120;
   assign soundFileAmplitudes [904] = 8'd127;
   assign soundFileAmplitudes [905] = 8'd123;
   assign soundFileAmplitudes [906] = 8'd120;
   assign soundFileAmplitudes [907] = 8'd116;
   assign soundFileAmplitudes [908] = 8'd129;
   assign soundFileAmplitudes [909] = 8'd140;
   assign soundFileAmplitudes [910] = 8'd149;
   assign soundFileAmplitudes [911] = 8'd148;
   assign soundFileAmplitudes [912] = 8'd133;
   assign soundFileAmplitudes [913] = 8'd113;
   assign soundFileAmplitudes [914] = 8'd103;
   assign soundFileAmplitudes [915] = 8'd113;
   assign soundFileAmplitudes [916] = 8'd121;
   assign soundFileAmplitudes [917] = 8'd107;
   assign soundFileAmplitudes [918] = 8'd92;
   assign soundFileAmplitudes [919] = 8'd103;
   assign soundFileAmplitudes [920] = 8'd118;
   assign soundFileAmplitudes [921] = 8'd129;
   assign soundFileAmplitudes [922] = 8'd126;
   assign soundFileAmplitudes [923] = 8'd129;
   assign soundFileAmplitudes [924] = 8'd137;
   assign soundFileAmplitudes [925] = 8'd148;
   assign soundFileAmplitudes [926] = 8'd153;
   assign soundFileAmplitudes [927] = 8'd145;
   assign soundFileAmplitudes [928] = 8'd143;
   assign soundFileAmplitudes [929] = 8'd139;
   assign soundFileAmplitudes [930] = 8'd141;
   assign soundFileAmplitudes [931] = 8'd148;
   assign soundFileAmplitudes [932] = 8'd138;
   assign soundFileAmplitudes [933] = 8'd120;
   assign soundFileAmplitudes [934] = 8'd117;
   assign soundFileAmplitudes [935] = 8'd128;
   assign soundFileAmplitudes [936] = 8'd135;
   assign soundFileAmplitudes [937] = 8'd135;
   assign soundFileAmplitudes [938] = 8'd133;
   assign soundFileAmplitudes [939] = 8'd124;
   assign soundFileAmplitudes [940] = 8'd117;
   assign soundFileAmplitudes [941] = 8'd116;
   assign soundFileAmplitudes [942] = 8'd131;
   assign soundFileAmplitudes [943] = 8'd133;
   assign soundFileAmplitudes [944] = 8'd126;
   assign soundFileAmplitudes [945] = 8'd124;
   assign soundFileAmplitudes [946] = 8'd122;
   assign soundFileAmplitudes [947] = 8'd111;
   assign soundFileAmplitudes [948] = 8'd79;
   assign soundFileAmplitudes [949] = 8'd87;
   assign soundFileAmplitudes [950] = 8'd101;
   assign soundFileAmplitudes [951] = 8'd110;
   assign soundFileAmplitudes [952] = 8'd114;
   assign soundFileAmplitudes [953] = 8'd112;
   assign soundFileAmplitudes [954] = 8'd125;
   assign soundFileAmplitudes [955] = 8'd133;
   assign soundFileAmplitudes [956] = 8'd146;
   assign soundFileAmplitudes [957] = 8'd145;
   assign soundFileAmplitudes [958] = 8'd145;
   assign soundFileAmplitudes [959] = 8'd155;
   assign soundFileAmplitudes [960] = 8'd153;
   assign soundFileAmplitudes [961] = 8'd148;
   assign soundFileAmplitudes [962] = 8'd149;
   assign soundFileAmplitudes [963] = 8'd154;
   assign soundFileAmplitudes [964] = 8'd143;
   assign soundFileAmplitudes [965] = 8'd133;
   assign soundFileAmplitudes [966] = 8'd134;
   assign soundFileAmplitudes [967] = 8'd128;
   assign soundFileAmplitudes [968] = 8'd122;
   assign soundFileAmplitudes [969] = 8'd118;
   assign soundFileAmplitudes [970] = 8'd126;
   assign soundFileAmplitudes [971] = 8'd129;
   assign soundFileAmplitudes [972] = 8'd126;
   assign soundFileAmplitudes [973] = 8'd123;
   assign soundFileAmplitudes [974] = 8'd118;
   assign soundFileAmplitudes [975] = 8'd116;
   assign soundFileAmplitudes [976] = 8'd108;
   assign soundFileAmplitudes [977] = 8'd106;
   assign soundFileAmplitudes [978] = 8'd102;
   assign soundFileAmplitudes [979] = 8'd107;
   assign soundFileAmplitudes [980] = 8'd115;
   assign soundFileAmplitudes [981] = 8'd119;
   assign soundFileAmplitudes [982] = 8'd108;
   assign soundFileAmplitudes [983] = 8'd89;
   assign soundFileAmplitudes [984] = 8'd101;
   assign soundFileAmplitudes [985] = 8'd116;
   assign soundFileAmplitudes [986] = 8'd124;
   assign soundFileAmplitudes [987] = 8'd136;
   assign soundFileAmplitudes [988] = 8'd137;
   assign soundFileAmplitudes [989] = 8'd128;
   assign soundFileAmplitudes [990] = 8'd136;
   assign soundFileAmplitudes [991] = 8'd142;
   assign soundFileAmplitudes [992] = 8'd144;
   assign soundFileAmplitudes [993] = 8'd151;
   assign soundFileAmplitudes [994] = 8'd150;
   assign soundFileAmplitudes [995] = 8'd138;
   assign soundFileAmplitudes [996] = 8'd135;
   assign soundFileAmplitudes [997] = 8'd140;
   assign soundFileAmplitudes [998] = 8'd134;
   assign soundFileAmplitudes [999] = 8'd136;
   assign soundFileAmplitudes [1000] = 8'd130;
   assign soundFileAmplitudes [1001] = 8'd126;
   assign soundFileAmplitudes [1002] = 8'd128;
   assign soundFileAmplitudes [1003] = 8'd117;
   assign soundFileAmplitudes [1004] = 8'd119;
   assign soundFileAmplitudes [1005] = 8'd131;
   assign soundFileAmplitudes [1006] = 8'd128;
   assign soundFileAmplitudes [1007] = 8'd118;
   assign soundFileAmplitudes [1008] = 8'd112;
   assign soundFileAmplitudes [1009] = 8'd113;
   assign soundFileAmplitudes [1010] = 8'd122;
   assign soundFileAmplitudes [1011] = 8'd128;
   assign soundFileAmplitudes [1012] = 8'd124;
   assign soundFileAmplitudes [1013] = 8'd120;
   assign soundFileAmplitudes [1014] = 8'd114;
   assign soundFileAmplitudes [1015] = 8'd129;
   assign soundFileAmplitudes [1016] = 8'd140;
   assign soundFileAmplitudes [1017] = 8'd138;
   assign soundFileAmplitudes [1018] = 8'd117;
   assign soundFileAmplitudes [1019] = 8'd107;
   assign soundFileAmplitudes [1020] = 8'd100;
   assign soundFileAmplitudes [1021] = 8'd105;
   assign soundFileAmplitudes [1022] = 8'd123;
   assign soundFileAmplitudes [1023] = 8'd123;
   assign soundFileAmplitudes [1024] = 8'd133;
   assign soundFileAmplitudes [1025] = 8'd116;
   assign soundFileAmplitudes [1026] = 8'd110;
   assign soundFileAmplitudes [1027] = 8'd119;
   assign soundFileAmplitudes [1028] = 8'd134;
   assign soundFileAmplitudes [1029] = 8'd146;
   assign soundFileAmplitudes [1030] = 8'd146;
   assign soundFileAmplitudes [1031] = 8'd139;
   assign soundFileAmplitudes [1032] = 8'd148;
   assign soundFileAmplitudes [1033] = 8'd147;
   assign soundFileAmplitudes [1034] = 8'd138;
   assign soundFileAmplitudes [1035] = 8'd141;
   assign soundFileAmplitudes [1036] = 8'd131;
   assign soundFileAmplitudes [1037] = 8'd122;
   assign soundFileAmplitudes [1038] = 8'd110;
   assign soundFileAmplitudes [1039] = 8'd109;
   assign soundFileAmplitudes [1040] = 8'd125;
   assign soundFileAmplitudes [1041] = 8'd135;
   assign soundFileAmplitudes [1042] = 8'd131;
   assign soundFileAmplitudes [1043] = 8'd122;
   assign soundFileAmplitudes [1044] = 8'd113;
   assign soundFileAmplitudes [1045] = 8'd118;
   assign soundFileAmplitudes [1046] = 8'd122;
   assign soundFileAmplitudes [1047] = 8'd132;
   assign soundFileAmplitudes [1048] = 8'd142;
   assign soundFileAmplitudes [1049] = 8'd137;
   assign soundFileAmplitudes [1050] = 8'd130;
   assign soundFileAmplitudes [1051] = 8'd138;
   assign soundFileAmplitudes [1052] = 8'd142;
   assign soundFileAmplitudes [1053] = 8'd127;
   assign soundFileAmplitudes [1054] = 8'd112;
   assign soundFileAmplitudes [1055] = 8'd98;
   assign soundFileAmplitudes [1056] = 8'd93;
   assign soundFileAmplitudes [1057] = 8'd98;
   assign soundFileAmplitudes [1058] = 8'd114;
   assign soundFileAmplitudes [1059] = 8'd121;
   assign soundFileAmplitudes [1060] = 8'd121;
   assign soundFileAmplitudes [1061] = 8'd121;
   assign soundFileAmplitudes [1062] = 8'd127;
   assign soundFileAmplitudes [1063] = 8'd144;
   assign soundFileAmplitudes [1064] = 8'd161;
   assign soundFileAmplitudes [1065] = 8'd153;
   assign soundFileAmplitudes [1066] = 8'd139;
   assign soundFileAmplitudes [1067] = 8'd143;
   assign soundFileAmplitudes [1068] = 8'd150;
   assign soundFileAmplitudes [1069] = 8'd148;
   assign soundFileAmplitudes [1070] = 8'd130;
   assign soundFileAmplitudes [1071] = 8'd126;
   assign soundFileAmplitudes [1072] = 8'd125;
   assign soundFileAmplitudes [1073] = 8'd123;
   assign soundFileAmplitudes [1074] = 8'd116;
   assign soundFileAmplitudes [1075] = 8'd109;
   assign soundFileAmplitudes [1076] = 8'd117;
   assign soundFileAmplitudes [1077] = 8'd125;
   assign soundFileAmplitudes [1078] = 8'd136;
   assign soundFileAmplitudes [1079] = 8'd139;
   assign soundFileAmplitudes [1080] = 8'd125;
   assign soundFileAmplitudes [1081] = 8'd126;
   assign soundFileAmplitudes [1082] = 8'd130;
   assign soundFileAmplitudes [1083] = 8'd132;
   assign soundFileAmplitudes [1084] = 8'd127;
   assign soundFileAmplitudes [1085] = 8'd128;
   assign soundFileAmplitudes [1086] = 8'd127;
   assign soundFileAmplitudes [1087] = 8'd110;
   assign soundFileAmplitudes [1088] = 8'd97;
   assign soundFileAmplitudes [1089] = 8'd99;
   assign soundFileAmplitudes [1090] = 8'd113;
   assign soundFileAmplitudes [1091] = 8'd120;
   assign soundFileAmplitudes [1092] = 8'd123;
   assign soundFileAmplitudes [1093] = 8'd122;
   assign soundFileAmplitudes [1094] = 8'd127;
   assign soundFileAmplitudes [1095] = 8'd118;
   assign soundFileAmplitudes [1096] = 8'd115;
   assign soundFileAmplitudes [1097] = 8'd119;
   assign soundFileAmplitudes [1098] = 8'd132;
   assign soundFileAmplitudes [1099] = 8'd153;
   assign soundFileAmplitudes [1100] = 8'd146;
   assign soundFileAmplitudes [1101] = 8'd125;
   assign soundFileAmplitudes [1102] = 8'd124;
   assign soundFileAmplitudes [1103] = 8'd128;
   assign soundFileAmplitudes [1104] = 8'd126;
   assign soundFileAmplitudes [1105] = 8'd125;
   assign soundFileAmplitudes [1106] = 8'd119;
   assign soundFileAmplitudes [1107] = 8'd119;
   assign soundFileAmplitudes [1108] = 8'd125;
   assign soundFileAmplitudes [1109] = 8'd143;
   assign soundFileAmplitudes [1110] = 8'd148;
   assign soundFileAmplitudes [1111] = 8'd147;
   assign soundFileAmplitudes [1112] = 8'd148;
   assign soundFileAmplitudes [1113] = 8'd139;
   assign soundFileAmplitudes [1114] = 8'd134;
   assign soundFileAmplitudes [1115] = 8'd128;
   assign soundFileAmplitudes [1116] = 8'd126;
   assign soundFileAmplitudes [1117] = 8'd124;
   assign soundFileAmplitudes [1118] = 8'd108;
   assign soundFileAmplitudes [1119] = 8'd101;
   assign soundFileAmplitudes [1120] = 8'd108;
   assign soundFileAmplitudes [1121] = 8'd120;
   assign soundFileAmplitudes [1122] = 8'd129;
   assign soundFileAmplitudes [1123] = 8'd113;
   assign soundFileAmplitudes [1124] = 8'd105;
   assign soundFileAmplitudes [1125] = 8'd116;
   assign soundFileAmplitudes [1126] = 8'd123;
   assign soundFileAmplitudes [1127] = 8'd122;
   assign soundFileAmplitudes [1128] = 8'd129;
   assign soundFileAmplitudes [1129] = 8'd136;
   assign soundFileAmplitudes [1130] = 8'd134;
   assign soundFileAmplitudes [1131] = 8'd126;
   assign soundFileAmplitudes [1132] = 8'd113;
   assign soundFileAmplitudes [1133] = 8'd121;
   assign soundFileAmplitudes [1134] = 8'd134;
   assign soundFileAmplitudes [1135] = 8'd133;
   assign soundFileAmplitudes [1136] = 8'd120;
   assign soundFileAmplitudes [1137] = 8'd115;
   assign soundFileAmplitudes [1138] = 8'd121;
   assign soundFileAmplitudes [1139] = 8'd126;
   assign soundFileAmplitudes [1140] = 8'd139;
   assign soundFileAmplitudes [1141] = 8'd144;
   assign soundFileAmplitudes [1142] = 8'd137;
   assign soundFileAmplitudes [1143] = 8'd140;
   assign soundFileAmplitudes [1144] = 8'd147;
   assign soundFileAmplitudes [1145] = 8'd147;
   assign soundFileAmplitudes [1146] = 8'd136;
   assign soundFileAmplitudes [1147] = 8'd142;
   assign soundFileAmplitudes [1148] = 8'd129;
   assign soundFileAmplitudes [1149] = 8'd111;
   assign soundFileAmplitudes [1150] = 8'd111;
   assign soundFileAmplitudes [1151] = 8'd114;
   assign soundFileAmplitudes [1152] = 8'd129;
   assign soundFileAmplitudes [1153] = 8'd128;
   assign soundFileAmplitudes [1154] = 8'd121;
   assign soundFileAmplitudes [1155] = 8'd119;
   assign soundFileAmplitudes [1156] = 8'd125;
   assign soundFileAmplitudes [1157] = 8'd140;
   assign soundFileAmplitudes [1158] = 8'd131;
   assign soundFileAmplitudes [1159] = 8'd102;
   assign soundFileAmplitudes [1160] = 8'd100;
   assign soundFileAmplitudes [1161] = 8'd114;
   assign soundFileAmplitudes [1162] = 8'd124;
   assign soundFileAmplitudes [1163] = 8'd108;
   assign soundFileAmplitudes [1164] = 8'd108;
   assign soundFileAmplitudes [1165] = 8'd101;
   assign soundFileAmplitudes [1166] = 8'd106;
   assign soundFileAmplitudes [1167] = 8'd116;
   assign soundFileAmplitudes [1168] = 8'd114;
   assign soundFileAmplitudes [1169] = 8'd129;
   assign soundFileAmplitudes [1170] = 8'd141;
   assign soundFileAmplitudes [1171] = 8'd146;
   assign soundFileAmplitudes [1172] = 8'd145;
   assign soundFileAmplitudes [1173] = 8'd149;
   assign soundFileAmplitudes [1174] = 8'd141;
   assign soundFileAmplitudes [1175] = 8'd144;
   assign soundFileAmplitudes [1176] = 8'd143;
   assign soundFileAmplitudes [1177] = 8'd139;
   assign soundFileAmplitudes [1178] = 8'd137;
   assign soundFileAmplitudes [1179] = 8'd129;
   assign soundFileAmplitudes [1180] = 8'd113;
   assign soundFileAmplitudes [1181] = 8'd110;
   assign soundFileAmplitudes [1182] = 8'd130;
   assign soundFileAmplitudes [1183] = 8'd143;
   assign soundFileAmplitudes [1184] = 8'd139;
   assign soundFileAmplitudes [1185] = 8'd133;
   assign soundFileAmplitudes [1186] = 8'd121;
   assign soundFileAmplitudes [1187] = 8'd124;
   assign soundFileAmplitudes [1188] = 8'd133;
   assign soundFileAmplitudes [1189] = 8'd133;
   assign soundFileAmplitudes [1190] = 8'd132;
   assign soundFileAmplitudes [1191] = 8'd134;
   assign soundFileAmplitudes [1192] = 8'd141;
   assign soundFileAmplitudes [1193] = 8'd129;
   assign soundFileAmplitudes [1194] = 8'd98;
   assign soundFileAmplitudes [1195] = 8'd90;
   assign soundFileAmplitudes [1196] = 8'd102;
   assign soundFileAmplitudes [1197] = 8'd102;
   assign soundFileAmplitudes [1198] = 8'd107;
   assign soundFileAmplitudes [1199] = 8'd103;
   assign soundFileAmplitudes [1200] = 8'd106;
   assign soundFileAmplitudes [1201] = 8'd111;
   assign soundFileAmplitudes [1202] = 8'd130;
   assign soundFileAmplitudes [1203] = 8'd146;
   assign soundFileAmplitudes [1204] = 8'd148;
   assign soundFileAmplitudes [1205] = 8'd151;
   assign soundFileAmplitudes [1206] = 8'd152;
   assign soundFileAmplitudes [1207] = 8'd151;
   assign soundFileAmplitudes [1208] = 8'd150;
   assign soundFileAmplitudes [1209] = 8'd151;
   assign soundFileAmplitudes [1210] = 8'd147;
   assign soundFileAmplitudes [1211] = 8'd126;
   assign soundFileAmplitudes [1212] = 8'd105;
   assign soundFileAmplitudes [1213] = 8'd110;
   assign soundFileAmplitudes [1214] = 8'd127;
   assign soundFileAmplitudes [1215] = 8'd136;
   assign soundFileAmplitudes [1216] = 8'd131;
   assign soundFileAmplitudes [1217] = 8'd124;
   assign soundFileAmplitudes [1218] = 8'd121;
   assign soundFileAmplitudes [1219] = 8'd122;
   assign soundFileAmplitudes [1220] = 8'd124;
   assign soundFileAmplitudes [1221] = 8'd126;
   assign soundFileAmplitudes [1222] = 8'd125;
   assign soundFileAmplitudes [1223] = 8'd135;
   assign soundFileAmplitudes [1224] = 8'd126;
   assign soundFileAmplitudes [1225] = 8'd111;
   assign soundFileAmplitudes [1226] = 8'd104;
   assign soundFileAmplitudes [1227] = 8'd110;
   assign soundFileAmplitudes [1228] = 8'd121;
   assign soundFileAmplitudes [1229] = 8'd119;
   assign soundFileAmplitudes [1230] = 8'd106;
   assign soundFileAmplitudes [1231] = 8'd99;
   assign soundFileAmplitudes [1232] = 8'd107;
   assign soundFileAmplitudes [1233] = 8'd116;
   assign soundFileAmplitudes [1234] = 8'd129;
   assign soundFileAmplitudes [1235] = 8'd135;
   assign soundFileAmplitudes [1236] = 8'd132;
   assign soundFileAmplitudes [1237] = 8'd139;
   assign soundFileAmplitudes [1238] = 8'd151;
   assign soundFileAmplitudes [1239] = 8'd151;
   assign soundFileAmplitudes [1240] = 8'd154;
   assign soundFileAmplitudes [1241] = 8'd151;
   assign soundFileAmplitudes [1242] = 8'd133;
   assign soundFileAmplitudes [1243] = 8'd124;
   assign soundFileAmplitudes [1244] = 8'd133;
   assign soundFileAmplitudes [1245] = 8'd137;
   assign soundFileAmplitudes [1246] = 8'd142;
   assign soundFileAmplitudes [1247] = 8'd138;
   assign soundFileAmplitudes [1248] = 8'd125;
   assign soundFileAmplitudes [1249] = 8'd118;
   assign soundFileAmplitudes [1250] = 8'd120;
   assign soundFileAmplitudes [1251] = 8'd120;
   assign soundFileAmplitudes [1252] = 8'd121;
   assign soundFileAmplitudes [1253] = 8'd115;
   assign soundFileAmplitudes [1254] = 8'd126;
   assign soundFileAmplitudes [1255] = 8'd133;
   assign soundFileAmplitudes [1256] = 8'd117;
   assign soundFileAmplitudes [1257] = 8'd107;
   assign soundFileAmplitudes [1258] = 8'd111;
   assign soundFileAmplitudes [1259] = 8'd116;
   assign soundFileAmplitudes [1260] = 8'd123;
   assign soundFileAmplitudes [1261] = 8'd123;
   assign soundFileAmplitudes [1262] = 8'd110;
   assign soundFileAmplitudes [1263] = 8'd112;
   assign soundFileAmplitudes [1264] = 8'd115;
   assign soundFileAmplitudes [1265] = 8'd132;
   assign soundFileAmplitudes [1266] = 8'd135;
   assign soundFileAmplitudes [1267] = 8'd121;
   assign soundFileAmplitudes [1268] = 8'd114;
   assign soundFileAmplitudes [1269] = 8'd129;
   assign soundFileAmplitudes [1270] = 8'd128;
   assign soundFileAmplitudes [1271] = 8'd128;
   assign soundFileAmplitudes [1272] = 8'd131;
   assign soundFileAmplitudes [1273] = 8'd128;
   assign soundFileAmplitudes [1274] = 8'd126;
   assign soundFileAmplitudes [1275] = 8'd124;
   assign soundFileAmplitudes [1276] = 8'd134;
   assign soundFileAmplitudes [1277] = 8'd146;
   assign soundFileAmplitudes [1278] = 8'd153;
   assign soundFileAmplitudes [1279] = 8'd144;
   assign soundFileAmplitudes [1280] = 8'd139;
   assign soundFileAmplitudes [1281] = 8'd140;
   assign soundFileAmplitudes [1282] = 8'd136;
   assign soundFileAmplitudes [1283] = 8'd129;
   assign soundFileAmplitudes [1284] = 8'd138;
   assign soundFileAmplitudes [1285] = 8'd135;
   assign soundFileAmplitudes [1286] = 8'd130;
   assign soundFileAmplitudes [1287] = 8'd108;
   assign soundFileAmplitudes [1288] = 8'd90;
   assign soundFileAmplitudes [1289] = 8'd100;
   assign soundFileAmplitudes [1290] = 8'd113;
   assign soundFileAmplitudes [1291] = 8'd120;
   assign soundFileAmplitudes [1292] = 8'd112;
   assign soundFileAmplitudes [1293] = 8'd107;
   assign soundFileAmplitudes [1294] = 8'd110;
   assign soundFileAmplitudes [1295] = 8'd114;
   assign soundFileAmplitudes [1296] = 8'd126;
   assign soundFileAmplitudes [1297] = 8'd134;
   assign soundFileAmplitudes [1298] = 8'd137;
   assign soundFileAmplitudes [1299] = 8'd133;
   assign soundFileAmplitudes [1300] = 8'd135;
   assign soundFileAmplitudes [1301] = 8'd141;
   assign soundFileAmplitudes [1302] = 8'd135;
   assign soundFileAmplitudes [1303] = 8'd129;
   assign soundFileAmplitudes [1304] = 8'd117;
   assign soundFileAmplitudes [1305] = 8'd101;
   assign soundFileAmplitudes [1306] = 8'd96;
   assign soundFileAmplitudes [1307] = 8'd107;
   assign soundFileAmplitudes [1308] = 8'd119;
   assign soundFileAmplitudes [1309] = 8'd130;
   assign soundFileAmplitudes [1310] = 8'd120;
   assign soundFileAmplitudes [1311] = 8'd123;
   assign soundFileAmplitudes [1312] = 8'd133;
   assign soundFileAmplitudes [1313] = 8'd154;
   assign soundFileAmplitudes [1314] = 8'd158;
   assign soundFileAmplitudes [1315] = 8'd158;
   assign soundFileAmplitudes [1316] = 8'd153;
   assign soundFileAmplitudes [1317] = 8'd153;
   assign soundFileAmplitudes [1318] = 8'd161;
   assign soundFileAmplitudes [1319] = 8'd143;
   assign soundFileAmplitudes [1320] = 8'd142;
   assign soundFileAmplitudes [1321] = 8'd129;
   assign soundFileAmplitudes [1322] = 8'd120;
   assign soundFileAmplitudes [1323] = 8'd112;
   assign soundFileAmplitudes [1324] = 8'd105;
   assign soundFileAmplitudes [1325] = 8'd99;
   assign soundFileAmplitudes [1326] = 8'd91;
   assign soundFileAmplitudes [1327] = 8'd97;
   assign soundFileAmplitudes [1328] = 8'd111;
   assign soundFileAmplitudes [1329] = 8'd117;
   assign soundFileAmplitudes [1330] = 8'd119;
   assign soundFileAmplitudes [1331] = 8'd116;
   assign soundFileAmplitudes [1332] = 8'd124;
   assign soundFileAmplitudes [1333] = 8'd141;
   assign soundFileAmplitudes [1334] = 8'd149;
   assign soundFileAmplitudes [1335] = 8'd146;
   assign soundFileAmplitudes [1336] = 8'd146;
   assign soundFileAmplitudes [1337] = 8'd143;
   assign soundFileAmplitudes [1338] = 8'd133;
   assign soundFileAmplitudes [1339] = 8'd117;
   assign soundFileAmplitudes [1340] = 8'd96;
   assign soundFileAmplitudes [1341] = 8'd99;
   assign soundFileAmplitudes [1342] = 8'd97;
   assign soundFileAmplitudes [1343] = 8'd114;
   assign soundFileAmplitudes [1344] = 8'd127;
   assign soundFileAmplitudes [1345] = 8'd125;
   assign soundFileAmplitudes [1346] = 8'd119;
   assign soundFileAmplitudes [1347] = 8'd119;
   assign soundFileAmplitudes [1348] = 8'd129;
   assign soundFileAmplitudes [1349] = 8'd161;
   assign soundFileAmplitudes [1350] = 8'd167;
   assign soundFileAmplitudes [1351] = 8'd149;
   assign soundFileAmplitudes [1352] = 8'd150;
   assign soundFileAmplitudes [1353] = 8'd148;
   assign soundFileAmplitudes [1354] = 8'd153;
   assign soundFileAmplitudes [1355] = 8'd142;
   assign soundFileAmplitudes [1356] = 8'd130;
   assign soundFileAmplitudes [1357] = 8'd122;
   assign soundFileAmplitudes [1358] = 8'd116;
   assign soundFileAmplitudes [1359] = 8'd115;
   assign soundFileAmplitudes [1360] = 8'd109;
   assign soundFileAmplitudes [1361] = 8'd112;
   assign soundFileAmplitudes [1362] = 8'd109;
   assign soundFileAmplitudes [1363] = 8'd112;
   assign soundFileAmplitudes [1364] = 8'd121;
   assign soundFileAmplitudes [1365] = 8'd114;
   assign soundFileAmplitudes [1366] = 8'd114;
   assign soundFileAmplitudes [1367] = 8'd119;
   assign soundFileAmplitudes [1368] = 8'd132;
   assign soundFileAmplitudes [1369] = 8'd132;
   assign soundFileAmplitudes [1370] = 8'd124;
   assign soundFileAmplitudes [1371] = 8'd124;
   assign soundFileAmplitudes [1372] = 8'd140;
   assign soundFileAmplitudes [1373] = 8'd148;
   assign soundFileAmplitudes [1374] = 8'd133;
   assign soundFileAmplitudes [1375] = 8'd102;
   assign soundFileAmplitudes [1376] = 8'd101;
   assign soundFileAmplitudes [1377] = 8'd114;
   assign soundFileAmplitudes [1378] = 8'd104;
   assign soundFileAmplitudes [1379] = 8'd115;
   assign soundFileAmplitudes [1380] = 8'd112;
   assign soundFileAmplitudes [1381] = 8'd118;
   assign soundFileAmplitudes [1382] = 8'd122;
   assign soundFileAmplitudes [1383] = 8'd116;
   assign soundFileAmplitudes [1384] = 8'd132;
   assign soundFileAmplitudes [1385] = 8'd155;
   assign soundFileAmplitudes [1386] = 8'd152;
   assign soundFileAmplitudes [1387] = 8'd141;
   assign soundFileAmplitudes [1388] = 8'd144;
   assign soundFileAmplitudes [1389] = 8'd141;
   assign soundFileAmplitudes [1390] = 8'd139;
   assign soundFileAmplitudes [1391] = 8'd142;
   assign soundFileAmplitudes [1392] = 8'd140;
   assign soundFileAmplitudes [1393] = 8'd134;
   assign soundFileAmplitudes [1394] = 8'd124;
   assign soundFileAmplitudes [1395] = 8'd121;
   assign soundFileAmplitudes [1396] = 8'd129;
   assign soundFileAmplitudes [1397] = 8'd127;
   assign soundFileAmplitudes [1398] = 8'd131;
   assign soundFileAmplitudes [1399] = 8'd126;
   assign soundFileAmplitudes [1400] = 8'd125;
   assign soundFileAmplitudes [1401] = 8'd108;
   assign soundFileAmplitudes [1402] = 8'd96;
   assign soundFileAmplitudes [1403] = 8'd114;
   assign soundFileAmplitudes [1404] = 8'd126;
   assign soundFileAmplitudes [1405] = 8'd124;
   assign soundFileAmplitudes [1406] = 8'd121;
   assign soundFileAmplitudes [1407] = 8'd127;
   assign soundFileAmplitudes [1408] = 8'd131;
   assign soundFileAmplitudes [1409] = 8'd120;
   assign soundFileAmplitudes [1410] = 8'd103;
   assign soundFileAmplitudes [1411] = 8'd107;
   assign soundFileAmplitudes [1412] = 8'd119;
   assign soundFileAmplitudes [1413] = 8'd119;
   assign soundFileAmplitudes [1414] = 8'd121;
   assign soundFileAmplitudes [1415] = 8'd125;
   assign soundFileAmplitudes [1416] = 8'd118;
   assign soundFileAmplitudes [1417] = 8'd112;
   assign soundFileAmplitudes [1418] = 8'd111;
   assign soundFileAmplitudes [1419] = 8'd114;
   assign soundFileAmplitudes [1420] = 8'd133;
   assign soundFileAmplitudes [1421] = 8'd145;
   assign soundFileAmplitudes [1422] = 8'd135;
   assign soundFileAmplitudes [1423] = 8'd137;
   assign soundFileAmplitudes [1424] = 8'd140;
   assign soundFileAmplitudes [1425] = 8'd148;
   assign soundFileAmplitudes [1426] = 8'd157;
   assign soundFileAmplitudes [1427] = 8'd151;
   assign soundFileAmplitudes [1428] = 8'd137;
   assign soundFileAmplitudes [1429] = 8'd134;
   assign soundFileAmplitudes [1430] = 8'd135;
   assign soundFileAmplitudes [1431] = 8'd134;
   assign soundFileAmplitudes [1432] = 8'd140;
   assign soundFileAmplitudes [1433] = 8'd137;
   assign soundFileAmplitudes [1434] = 8'd128;
   assign soundFileAmplitudes [1435] = 8'd114;
   assign soundFileAmplitudes [1436] = 8'd112;
   assign soundFileAmplitudes [1437] = 8'd114;
   assign soundFileAmplitudes [1438] = 8'd117;
   assign soundFileAmplitudes [1439] = 8'd123;
   assign soundFileAmplitudes [1440] = 8'd119;
   assign soundFileAmplitudes [1441] = 8'd118;
   assign soundFileAmplitudes [1442] = 8'd120;
   assign soundFileAmplitudes [1443] = 8'd122;
   assign soundFileAmplitudes [1444] = 8'd119;
   assign soundFileAmplitudes [1445] = 8'd102;
   assign soundFileAmplitudes [1446] = 8'd107;
   assign soundFileAmplitudes [1447] = 8'd122;
   assign soundFileAmplitudes [1448] = 8'd117;
   assign soundFileAmplitudes [1449] = 8'd116;
   assign soundFileAmplitudes [1450] = 8'd113;
   assign soundFileAmplitudes [1451] = 8'd113;
   assign soundFileAmplitudes [1452] = 8'd113;
   assign soundFileAmplitudes [1453] = 8'd119;
   assign soundFileAmplitudes [1454] = 8'd120;
   assign soundFileAmplitudes [1455] = 8'd131;
   assign soundFileAmplitudes [1456] = 8'd145;
   assign soundFileAmplitudes [1457] = 8'd141;
   assign soundFileAmplitudes [1458] = 8'd148;
   assign soundFileAmplitudes [1459] = 8'd154;
   assign soundFileAmplitudes [1460] = 8'd148;
   assign soundFileAmplitudes [1461] = 8'd148;
   assign soundFileAmplitudes [1462] = 8'd149;
   assign soundFileAmplitudes [1463] = 8'd137;
   assign soundFileAmplitudes [1464] = 8'd133;
   assign soundFileAmplitudes [1465] = 8'd128;
   assign soundFileAmplitudes [1466] = 8'd124;
   assign soundFileAmplitudes [1467] = 8'd119;
   assign soundFileAmplitudes [1468] = 8'd130;
   assign soundFileAmplitudes [1469] = 8'd131;
   assign soundFileAmplitudes [1470] = 8'd129;
   assign soundFileAmplitudes [1471] = 8'd121;
   assign soundFileAmplitudes [1472] = 8'd111;
   assign soundFileAmplitudes [1473] = 8'd118;
   assign soundFileAmplitudes [1474] = 8'd121;
   assign soundFileAmplitudes [1475] = 8'd122;
   assign soundFileAmplitudes [1476] = 8'd114;
   assign soundFileAmplitudes [1477] = 8'd116;
   assign soundFileAmplitudes [1478] = 8'd126;
   assign soundFileAmplitudes [1479] = 8'd131;
   assign soundFileAmplitudes [1480] = 8'd115;
   assign soundFileAmplitudes [1481] = 8'd113;
   assign soundFileAmplitudes [1482] = 8'd121;
   assign soundFileAmplitudes [1483] = 8'd119;
   assign soundFileAmplitudes [1484] = 8'd112;
   assign soundFileAmplitudes [1485] = 8'd109;
   assign soundFileAmplitudes [1486] = 8'd109;
   assign soundFileAmplitudes [1487] = 8'd116;
   assign soundFileAmplitudes [1488] = 8'd131;
   assign soundFileAmplitudes [1489] = 8'd138;
   assign soundFileAmplitudes [1490] = 8'd144;
   assign soundFileAmplitudes [1491] = 8'd158;
   assign soundFileAmplitudes [1492] = 8'd161;
   assign soundFileAmplitudes [1493] = 8'd151;
   assign soundFileAmplitudes [1494] = 8'd153;
   assign soundFileAmplitudes [1495] = 8'd144;
   assign soundFileAmplitudes [1496] = 8'd139;
   assign soundFileAmplitudes [1497] = 8'd140;
   assign soundFileAmplitudes [1498] = 8'd132;
   assign soundFileAmplitudes [1499] = 8'd126;
   assign soundFileAmplitudes [1500] = 8'd116;
   assign soundFileAmplitudes [1501] = 8'd112;
   assign soundFileAmplitudes [1502] = 8'd119;
   assign soundFileAmplitudes [1503] = 8'd120;
   assign soundFileAmplitudes [1504] = 8'd117;
   assign soundFileAmplitudes [1505] = 8'd121;
   assign soundFileAmplitudes [1506] = 8'd112;
   assign soundFileAmplitudes [1507] = 8'd113;
   assign soundFileAmplitudes [1508] = 8'd112;
   assign soundFileAmplitudes [1509] = 8'd118;
   assign soundFileAmplitudes [1510] = 8'd125;
   assign soundFileAmplitudes [1511] = 8'd119;
   assign soundFileAmplitudes [1512] = 8'd126;
   assign soundFileAmplitudes [1513] = 8'd129;
   assign soundFileAmplitudes [1514] = 8'd125;
   assign soundFileAmplitudes [1515] = 8'd97;
   assign soundFileAmplitudes [1516] = 8'd93;
   assign soundFileAmplitudes [1517] = 8'd101;
   assign soundFileAmplitudes [1518] = 8'd112;
   assign soundFileAmplitudes [1519] = 8'd118;
   assign soundFileAmplitudes [1520] = 8'd116;
   assign soundFileAmplitudes [1521] = 8'd120;
   assign soundFileAmplitudes [1522] = 8'd114;
   assign soundFileAmplitudes [1523] = 8'd128;
   assign soundFileAmplitudes [1524] = 8'd135;
   assign soundFileAmplitudes [1525] = 8'd152;
   assign soundFileAmplitudes [1526] = 8'd168;
   assign soundFileAmplitudes [1527] = 8'd174;
   assign soundFileAmplitudes [1528] = 8'd165;
   assign soundFileAmplitudes [1529] = 8'd157;
   assign soundFileAmplitudes [1530] = 8'd158;
   assign soundFileAmplitudes [1531] = 8'd141;
   assign soundFileAmplitudes [1532] = 8'd133;
   assign soundFileAmplitudes [1533] = 8'd125;
   assign soundFileAmplitudes [1534] = 8'd120;
   assign soundFileAmplitudes [1535] = 8'd113;
   assign soundFileAmplitudes [1536] = 8'd108;
   assign soundFileAmplitudes [1537] = 8'd109;
   assign soundFileAmplitudes [1538] = 8'd111;
   assign soundFileAmplitudes [1539] = 8'd115;
   assign soundFileAmplitudes [1540] = 8'd112;
   assign soundFileAmplitudes [1541] = 8'd116;
   assign soundFileAmplitudes [1542] = 8'd121;
   assign soundFileAmplitudes [1543] = 8'd124;
   assign soundFileAmplitudes [1544] = 8'd126;
   assign soundFileAmplitudes [1545] = 8'd124;
   assign soundFileAmplitudes [1546] = 8'd120;
   assign soundFileAmplitudes [1547] = 8'd124;
   assign soundFileAmplitudes [1548] = 8'd128;
   assign soundFileAmplitudes [1549] = 8'd106;
   assign soundFileAmplitudes [1550] = 8'd104;
   assign soundFileAmplitudes [1551] = 8'd107;
   assign soundFileAmplitudes [1552] = 8'd104;
   assign soundFileAmplitudes [1553] = 8'd109;
   assign soundFileAmplitudes [1554] = 8'd108;
   assign soundFileAmplitudes [1555] = 8'd111;
   assign soundFileAmplitudes [1556] = 8'd124;
   assign soundFileAmplitudes [1557] = 8'd132;
   assign soundFileAmplitudes [1558] = 8'd137;
   assign soundFileAmplitudes [1559] = 8'd152;
   assign soundFileAmplitudes [1560] = 8'd156;
   assign soundFileAmplitudes [1561] = 8'd167;
   assign soundFileAmplitudes [1562] = 8'd163;
   assign soundFileAmplitudes [1563] = 8'd159;
   assign soundFileAmplitudes [1564] = 8'd160;
   assign soundFileAmplitudes [1565] = 8'd161;
   assign soundFileAmplitudes [1566] = 8'd157;
   assign soundFileAmplitudes [1567] = 8'd142;
   assign soundFileAmplitudes [1568] = 8'd129;
   assign soundFileAmplitudes [1569] = 8'd112;
   assign soundFileAmplitudes [1570] = 8'd98;
   assign soundFileAmplitudes [1571] = 8'd95;
   assign soundFileAmplitudes [1572] = 8'd103;
   assign soundFileAmplitudes [1573] = 8'd115;
   assign soundFileAmplitudes [1574] = 8'd113;
   assign soundFileAmplitudes [1575] = 8'd97;
   assign soundFileAmplitudes [1576] = 8'd103;
   assign soundFileAmplitudes [1577] = 8'd108;
   assign soundFileAmplitudes [1578] = 8'd118;
   assign soundFileAmplitudes [1579] = 8'd129;
   assign soundFileAmplitudes [1580] = 8'd135;
   assign soundFileAmplitudes [1581] = 8'd125;
   assign soundFileAmplitudes [1582] = 8'd131;
   assign soundFileAmplitudes [1583] = 8'd122;
   assign soundFileAmplitudes [1584] = 8'd106;
   assign soundFileAmplitudes [1585] = 8'd120;
   assign soundFileAmplitudes [1586] = 8'd111;
   assign soundFileAmplitudes [1587] = 8'd110;
   assign soundFileAmplitudes [1588] = 8'd113;
   assign soundFileAmplitudes [1589] = 8'd116;
   assign soundFileAmplitudes [1590] = 8'd124;
   assign soundFileAmplitudes [1591] = 8'd137;
   assign soundFileAmplitudes [1592] = 8'd132;
   assign soundFileAmplitudes [1593] = 8'd131;
   assign soundFileAmplitudes [1594] = 8'd131;
   assign soundFileAmplitudes [1595] = 8'd137;
   assign soundFileAmplitudes [1596] = 8'd156;
   assign soundFileAmplitudes [1597] = 8'd165;
   assign soundFileAmplitudes [1598] = 8'd161;
   assign soundFileAmplitudes [1599] = 8'd156;
   assign soundFileAmplitudes [1600] = 8'd150;
   assign soundFileAmplitudes [1601] = 8'd140;
   assign soundFileAmplitudes [1602] = 8'd143;
   assign soundFileAmplitudes [1603] = 8'd135;
   assign soundFileAmplitudes [1604] = 8'd129;
   assign soundFileAmplitudes [1605] = 8'd116;
   assign soundFileAmplitudes [1606] = 8'd108;
   assign soundFileAmplitudes [1607] = 8'd113;
   assign soundFileAmplitudes [1608] = 8'd111;
   assign soundFileAmplitudes [1609] = 8'd103;
   assign soundFileAmplitudes [1610] = 8'd101;
   assign soundFileAmplitudes [1611] = 8'd101;
   assign soundFileAmplitudes [1612] = 8'd115;
   assign soundFileAmplitudes [1613] = 8'd125;
   assign soundFileAmplitudes [1614] = 8'd137;
   assign soundFileAmplitudes [1615] = 8'd133;
   assign soundFileAmplitudes [1616] = 8'd120;
   assign soundFileAmplitudes [1617] = 8'd128;
   assign soundFileAmplitudes [1618] = 8'd114;
   assign soundFileAmplitudes [1619] = 8'd112;
   assign soundFileAmplitudes [1620] = 8'd119;
   assign soundFileAmplitudes [1621] = 8'd122;
   assign soundFileAmplitudes [1622] = 8'd119;
   assign soundFileAmplitudes [1623] = 8'd125;
   assign soundFileAmplitudes [1624] = 8'd118;
   assign soundFileAmplitudes [1625] = 8'd125;
   assign soundFileAmplitudes [1626] = 8'd133;
   assign soundFileAmplitudes [1627] = 8'd124;
   assign soundFileAmplitudes [1628] = 8'd139;
   assign soundFileAmplitudes [1629] = 8'd138;
   assign soundFileAmplitudes [1630] = 8'd139;
   assign soundFileAmplitudes [1631] = 8'd147;
   assign soundFileAmplitudes [1632] = 8'd147;
   assign soundFileAmplitudes [1633] = 8'd144;
   assign soundFileAmplitudes [1634] = 8'd142;
   assign soundFileAmplitudes [1635] = 8'd138;
   assign soundFileAmplitudes [1636] = 8'd141;
   assign soundFileAmplitudes [1637] = 8'd136;
   assign soundFileAmplitudes [1638] = 8'd130;
   assign soundFileAmplitudes [1639] = 8'd119;
   assign soundFileAmplitudes [1640] = 8'd111;
   assign soundFileAmplitudes [1641] = 8'd106;
   assign soundFileAmplitudes [1642] = 8'd110;
   assign soundFileAmplitudes [1643] = 8'd115;
   assign soundFileAmplitudes [1644] = 8'd114;
   assign soundFileAmplitudes [1645] = 8'd114;
   assign soundFileAmplitudes [1646] = 8'd105;
   assign soundFileAmplitudes [1647] = 8'd113;
   assign soundFileAmplitudes [1648] = 8'd119;
   assign soundFileAmplitudes [1649] = 8'd135;
   assign soundFileAmplitudes [1650] = 8'd131;
   assign soundFileAmplitudes [1651] = 8'd133;
   assign soundFileAmplitudes [1652] = 8'd129;
   assign soundFileAmplitudes [1653] = 8'd108;
   assign soundFileAmplitudes [1654] = 8'd111;
   assign soundFileAmplitudes [1655] = 8'd114;
   assign soundFileAmplitudes [1656] = 8'd115;
   assign soundFileAmplitudes [1657] = 8'd116;
   assign soundFileAmplitudes [1658] = 8'd127;
   assign soundFileAmplitudes [1659] = 8'd130;
   assign soundFileAmplitudes [1660] = 8'd139;
   assign soundFileAmplitudes [1661] = 8'd134;
   assign soundFileAmplitudes [1662] = 8'd137;
   assign soundFileAmplitudes [1663] = 8'd141;
   assign soundFileAmplitudes [1664] = 8'd140;
   assign soundFileAmplitudes [1665] = 8'd152;
   assign soundFileAmplitudes [1666] = 8'd152;
   assign soundFileAmplitudes [1667] = 8'd150;
   assign soundFileAmplitudes [1668] = 8'd139;
   assign soundFileAmplitudes [1669] = 8'd131;
   assign soundFileAmplitudes [1670] = 8'd127;
   assign soundFileAmplitudes [1671] = 8'd126;
   assign soundFileAmplitudes [1672] = 8'd117;
   assign soundFileAmplitudes [1673] = 8'd110;
   assign soundFileAmplitudes [1674] = 8'd106;
   assign soundFileAmplitudes [1675] = 8'd110;
   assign soundFileAmplitudes [1676] = 8'd112;
   assign soundFileAmplitudes [1677] = 8'd120;
   assign soundFileAmplitudes [1678] = 8'd120;
   assign soundFileAmplitudes [1679] = 8'd113;
   assign soundFileAmplitudes [1680] = 8'd115;
   assign soundFileAmplitudes [1681] = 8'd119;
   assign soundFileAmplitudes [1682] = 8'd131;
   assign soundFileAmplitudes [1683] = 8'd142;
   assign soundFileAmplitudes [1684] = 8'd141;
   assign soundFileAmplitudes [1685] = 8'd130;
   assign soundFileAmplitudes [1686] = 8'd130;
   assign soundFileAmplitudes [1687] = 8'd109;
   assign soundFileAmplitudes [1688] = 8'd105;
   assign soundFileAmplitudes [1689] = 8'd111;
   assign soundFileAmplitudes [1690] = 8'd113;
   assign soundFileAmplitudes [1691] = 8'd118;
   assign soundFileAmplitudes [1692] = 8'd121;
   assign soundFileAmplitudes [1693] = 8'd119;
   assign soundFileAmplitudes [1694] = 8'd129;
   assign soundFileAmplitudes [1695] = 8'd138;
   assign soundFileAmplitudes [1696] = 8'd133;
   assign soundFileAmplitudes [1697] = 8'd139;
   assign soundFileAmplitudes [1698] = 8'd132;
   assign soundFileAmplitudes [1699] = 8'd142;
   assign soundFileAmplitudes [1700] = 8'd154;
   assign soundFileAmplitudes [1701] = 8'd157;
   assign soundFileAmplitudes [1702] = 8'd147;
   assign soundFileAmplitudes [1703] = 8'd137;
   assign soundFileAmplitudes [1704] = 8'd126;
   assign soundFileAmplitudes [1705] = 8'd125;
   assign soundFileAmplitudes [1706] = 8'd125;
   assign soundFileAmplitudes [1707] = 8'd121;
   assign soundFileAmplitudes [1708] = 8'd110;
   assign soundFileAmplitudes [1709] = 8'd102;
   assign soundFileAmplitudes [1710] = 8'd104;
   assign soundFileAmplitudes [1711] = 8'd102;
   assign soundFileAmplitudes [1712] = 8'd111;
   assign soundFileAmplitudes [1713] = 8'd111;
   assign soundFileAmplitudes [1714] = 8'd114;
   assign soundFileAmplitudes [1715] = 8'd111;
   assign soundFileAmplitudes [1716] = 8'd121;
   assign soundFileAmplitudes [1717] = 8'd131;
   assign soundFileAmplitudes [1718] = 8'd133;
   assign soundFileAmplitudes [1719] = 8'd137;
   assign soundFileAmplitudes [1720] = 8'd141;
   assign soundFileAmplitudes [1721] = 8'd141;
   assign soundFileAmplitudes [1722] = 8'd128;
   assign soundFileAmplitudes [1723] = 8'd127;
   assign soundFileAmplitudes [1724] = 8'd137;
   assign soundFileAmplitudes [1725] = 8'd136;
   assign soundFileAmplitudes [1726] = 8'd131;
   assign soundFileAmplitudes [1727] = 8'd124;
   assign soundFileAmplitudes [1728] = 8'd116;
   assign soundFileAmplitudes [1729] = 8'd132;
   assign soundFileAmplitudes [1730] = 8'd127;
   assign soundFileAmplitudes [1731] = 8'd130;
   assign soundFileAmplitudes [1732] = 8'd134;
   assign soundFileAmplitudes [1733] = 8'd135;
   assign soundFileAmplitudes [1734] = 8'd150;
   assign soundFileAmplitudes [1735] = 8'd148;
   assign soundFileAmplitudes [1736] = 8'd138;
   assign soundFileAmplitudes [1737] = 8'd132;
   assign soundFileAmplitudes [1738] = 8'd139;
   assign soundFileAmplitudes [1739] = 8'd142;
   assign soundFileAmplitudes [1740] = 8'd138;
   assign soundFileAmplitudes [1741] = 8'd123;
   assign soundFileAmplitudes [1742] = 8'd108;
   assign soundFileAmplitudes [1743] = 8'd103;
   assign soundFileAmplitudes [1744] = 8'd103;
   assign soundFileAmplitudes [1745] = 8'd104;
   assign soundFileAmplitudes [1746] = 8'd113;
   assign soundFileAmplitudes [1747] = 8'd115;
   assign soundFileAmplitudes [1748] = 8'd113;
   assign soundFileAmplitudes [1749] = 8'd108;
   assign soundFileAmplitudes [1750] = 8'd103;
   assign soundFileAmplitudes [1751] = 8'd112;
   assign soundFileAmplitudes [1752] = 8'd118;
   assign soundFileAmplitudes [1753] = 8'd132;
   assign soundFileAmplitudes [1754] = 8'd138;
   assign soundFileAmplitudes [1755] = 8'd139;
   assign soundFileAmplitudes [1756] = 8'd131;
   assign soundFileAmplitudes [1757] = 8'd114;
   assign soundFileAmplitudes [1758] = 8'd125;
   assign soundFileAmplitudes [1759] = 8'd136;
   assign soundFileAmplitudes [1760] = 8'd134;
   assign soundFileAmplitudes [1761] = 8'd132;
   assign soundFileAmplitudes [1762] = 8'd121;
   assign soundFileAmplitudes [1763] = 8'd129;
   assign soundFileAmplitudes [1764] = 8'd130;
   assign soundFileAmplitudes [1765] = 8'd127;
   assign soundFileAmplitudes [1766] = 8'd128;
   assign soundFileAmplitudes [1767] = 8'd127;
   assign soundFileAmplitudes [1768] = 8'd143;
   assign soundFileAmplitudes [1769] = 8'd152;
   assign soundFileAmplitudes [1770] = 8'd146;
   assign soundFileAmplitudes [1771] = 8'd134;
   assign soundFileAmplitudes [1772] = 8'd128;
   assign soundFileAmplitudes [1773] = 8'd132;
   assign soundFileAmplitudes [1774] = 8'd137;
   assign soundFileAmplitudes [1775] = 8'd129;
   assign soundFileAmplitudes [1776] = 8'd112;
   assign soundFileAmplitudes [1777] = 8'd101;
   assign soundFileAmplitudes [1778] = 8'd102;
   assign soundFileAmplitudes [1779] = 8'd116;
   assign soundFileAmplitudes [1780] = 8'd127;
   assign soundFileAmplitudes [1781] = 8'd132;
   assign soundFileAmplitudes [1782] = 8'd126;
   assign soundFileAmplitudes [1783] = 8'd124;
   assign soundFileAmplitudes [1784] = 8'd122;
   assign soundFileAmplitudes [1785] = 8'd125;
   assign soundFileAmplitudes [1786] = 8'd138;
   assign soundFileAmplitudes [1787] = 8'd137;
   assign soundFileAmplitudes [1788] = 8'd137;
   assign soundFileAmplitudes [1789] = 8'd136;
   assign soundFileAmplitudes [1790] = 8'd132;
   assign soundFileAmplitudes [1791] = 8'd113;
   assign soundFileAmplitudes [1792] = 8'd104;
   assign soundFileAmplitudes [1793] = 8'd115;
   assign soundFileAmplitudes [1794] = 8'd114;
   assign soundFileAmplitudes [1795] = 8'd116;
   assign soundFileAmplitudes [1796] = 8'd119;
   assign soundFileAmplitudes [1797] = 8'd120;
   assign soundFileAmplitudes [1798] = 8'd128;
   assign soundFileAmplitudes [1799] = 8'd123;
   assign soundFileAmplitudes [1800] = 8'd130;
   assign soundFileAmplitudes [1801] = 8'd143;
   assign soundFileAmplitudes [1802] = 8'd150;
   assign soundFileAmplitudes [1803] = 8'd164;
   assign soundFileAmplitudes [1804] = 8'd153;
   assign soundFileAmplitudes [1805] = 8'd144;
   assign soundFileAmplitudes [1806] = 8'd141;
   assign soundFileAmplitudes [1807] = 8'd129;
   assign soundFileAmplitudes [1808] = 8'd121;
   assign soundFileAmplitudes [1809] = 8'd116;
   assign soundFileAmplitudes [1810] = 8'd102;
   assign soundFileAmplitudes [1811] = 8'd95;
   assign soundFileAmplitudes [1812] = 8'd91;
   assign soundFileAmplitudes [1813] = 8'd91;
   assign soundFileAmplitudes [1814] = 8'd99;
   assign soundFileAmplitudes [1815] = 8'd105;
   assign soundFileAmplitudes [1816] = 8'd114;
   assign soundFileAmplitudes [1817] = 8'd117;
   assign soundFileAmplitudes [1818] = 8'd128;
   assign soundFileAmplitudes [1819] = 8'd137;
   assign soundFileAmplitudes [1820] = 8'd144;
   assign soundFileAmplitudes [1821] = 8'd152;
   assign soundFileAmplitudes [1822] = 8'd149;
   assign soundFileAmplitudes [1823] = 8'd144;
   assign soundFileAmplitudes [1824] = 8'd145;
   assign soundFileAmplitudes [1825] = 8'd130;
   assign soundFileAmplitudes [1826] = 8'd118;
   assign soundFileAmplitudes [1827] = 8'd119;
   assign soundFileAmplitudes [1828] = 8'd110;
   assign soundFileAmplitudes [1829] = 8'd104;
   assign soundFileAmplitudes [1830] = 8'd105;
   assign soundFileAmplitudes [1831] = 8'd106;
   assign soundFileAmplitudes [1832] = 8'd122;
   assign soundFileAmplitudes [1833] = 8'd125;
   assign soundFileAmplitudes [1834] = 8'd124;
   assign soundFileAmplitudes [1835] = 8'd138;
   assign soundFileAmplitudes [1836] = 8'd142;
   assign soundFileAmplitudes [1837] = 8'd149;
   assign soundFileAmplitudes [1838] = 8'd160;
   assign soundFileAmplitudes [1839] = 8'd153;
   assign soundFileAmplitudes [1840] = 8'd152;
   assign soundFileAmplitudes [1841] = 8'd150;
   assign soundFileAmplitudes [1842] = 8'd152;
   assign soundFileAmplitudes [1843] = 8'd153;
   assign soundFileAmplitudes [1844] = 8'd121;
   assign soundFileAmplitudes [1845] = 8'd98;
   assign soundFileAmplitudes [1846] = 8'd81;
   assign soundFileAmplitudes [1847] = 8'd88;
   assign soundFileAmplitudes [1848] = 8'd99;
   assign soundFileAmplitudes [1849] = 8'd103;
   assign soundFileAmplitudes [1850] = 8'd106;
   assign soundFileAmplitudes [1851] = 8'd105;
   assign soundFileAmplitudes [1852] = 8'd107;
   assign soundFileAmplitudes [1853] = 8'd107;
   assign soundFileAmplitudes [1854] = 8'd120;
   assign soundFileAmplitudes [1855] = 8'd137;
   assign soundFileAmplitudes [1856] = 8'd152;
   assign soundFileAmplitudes [1857] = 8'd153;
   assign soundFileAmplitudes [1858] = 8'd158;
   assign soundFileAmplitudes [1859] = 8'd155;
   assign soundFileAmplitudes [1860] = 8'd143;
   assign soundFileAmplitudes [1861] = 8'd135;
   assign soundFileAmplitudes [1862] = 8'd130;
   assign soundFileAmplitudes [1863] = 8'd119;
   assign soundFileAmplitudes [1864] = 8'd115;
   assign soundFileAmplitudes [1865] = 8'd119;
   assign soundFileAmplitudes [1866] = 8'd118;
   assign soundFileAmplitudes [1867] = 8'd113;
   assign soundFileAmplitudes [1868] = 8'd105;
   assign soundFileAmplitudes [1869] = 8'd114;
   assign soundFileAmplitudes [1870] = 8'd129;
   assign soundFileAmplitudes [1871] = 8'd138;
   assign soundFileAmplitudes [1872] = 8'd148;
   assign soundFileAmplitudes [1873] = 8'd153;
   assign soundFileAmplitudes [1874] = 8'd148;
   assign soundFileAmplitudes [1875] = 8'd148;
   assign soundFileAmplitudes [1876] = 8'd152;
   assign soundFileAmplitudes [1877] = 8'd136;
   assign soundFileAmplitudes [1878] = 8'd126;
   assign soundFileAmplitudes [1879] = 8'd129;
   assign soundFileAmplitudes [1880] = 8'd112;
   assign soundFileAmplitudes [1881] = 8'd109;
   assign soundFileAmplitudes [1882] = 8'd106;
   assign soundFileAmplitudes [1883] = 8'd104;
   assign soundFileAmplitudes [1884] = 8'd111;
   assign soundFileAmplitudes [1885] = 8'd103;
   assign soundFileAmplitudes [1886] = 8'd99;
   assign soundFileAmplitudes [1887] = 8'd100;
   assign soundFileAmplitudes [1888] = 8'd109;
   assign soundFileAmplitudes [1889] = 8'd116;
   assign soundFileAmplitudes [1890] = 8'd120;
   assign soundFileAmplitudes [1891] = 8'd131;
   assign soundFileAmplitudes [1892] = 8'd142;
   assign soundFileAmplitudes [1893] = 8'd150;
   assign soundFileAmplitudes [1894] = 8'd142;
   assign soundFileAmplitudes [1895] = 8'd135;
   assign soundFileAmplitudes [1896] = 8'd136;
   assign soundFileAmplitudes [1897] = 8'd138;
   assign soundFileAmplitudes [1898] = 8'd132;
   assign soundFileAmplitudes [1899] = 8'd124;
   assign soundFileAmplitudes [1900] = 8'd120;
   assign soundFileAmplitudes [1901] = 8'd120;
   assign soundFileAmplitudes [1902] = 8'd134;
   assign soundFileAmplitudes [1903] = 8'd140;
   assign soundFileAmplitudes [1904] = 8'd139;
   assign soundFileAmplitudes [1905] = 8'd131;
   assign soundFileAmplitudes [1906] = 8'd133;
   assign soundFileAmplitudes [1907] = 8'd141;
   assign soundFileAmplitudes [1908] = 8'd148;
   assign soundFileAmplitudes [1909] = 8'd136;
   assign soundFileAmplitudes [1910] = 8'd131;
   assign soundFileAmplitudes [1911] = 8'd128;
   assign soundFileAmplitudes [1912] = 8'd123;
   assign soundFileAmplitudes [1913] = 8'd122;
   assign soundFileAmplitudes [1914] = 8'd113;
   assign soundFileAmplitudes [1915] = 8'd117;
   assign soundFileAmplitudes [1916] = 8'd112;
   assign soundFileAmplitudes [1917] = 8'd112;
   assign soundFileAmplitudes [1918] = 8'd111;
   assign soundFileAmplitudes [1919] = 8'd107;
   assign soundFileAmplitudes [1920] = 8'd115;
   assign soundFileAmplitudes [1921] = 8'd120;
   assign soundFileAmplitudes [1922] = 8'd116;
   assign soundFileAmplitudes [1923] = 8'd120;
   assign soundFileAmplitudes [1924] = 8'd111;
   assign soundFileAmplitudes [1925] = 8'd110;
   assign soundFileAmplitudes [1926] = 8'd116;
   assign soundFileAmplitudes [1927] = 8'd122;
   assign soundFileAmplitudes [1928] = 8'd138;
   assign soundFileAmplitudes [1929] = 8'd137;
   assign soundFileAmplitudes [1930] = 8'd130;
   assign soundFileAmplitudes [1931] = 8'd131;
   assign soundFileAmplitudes [1932] = 8'd132;
   assign soundFileAmplitudes [1933] = 8'd129;
   assign soundFileAmplitudes [1934] = 8'd130;
   assign soundFileAmplitudes [1935] = 8'd135;
   assign soundFileAmplitudes [1936] = 8'd142;
   assign soundFileAmplitudes [1937] = 8'd142;
   assign soundFileAmplitudes [1938] = 8'd134;
   assign soundFileAmplitudes [1939] = 8'd137;
   assign soundFileAmplitudes [1940] = 8'd137;
   assign soundFileAmplitudes [1941] = 8'd133;
   assign soundFileAmplitudes [1942] = 8'd142;
   assign soundFileAmplitudes [1943] = 8'd139;
   assign soundFileAmplitudes [1944] = 8'd141;
   assign soundFileAmplitudes [1945] = 8'd137;
   assign soundFileAmplitudes [1946] = 8'd125;
   assign soundFileAmplitudes [1947] = 8'd118;
   assign soundFileAmplitudes [1948] = 8'd109;
   assign soundFileAmplitudes [1949] = 8'd106;
   assign soundFileAmplitudes [1950] = 8'd107;
   assign soundFileAmplitudes [1951] = 8'd119;
   assign soundFileAmplitudes [1952] = 8'd121;
   assign soundFileAmplitudes [1953] = 8'd118;
   assign soundFileAmplitudes [1954] = 8'd115;
   assign soundFileAmplitudes [1955] = 8'd113;
   assign soundFileAmplitudes [1956] = 8'd117;
   assign soundFileAmplitudes [1957] = 8'd123;
   assign soundFileAmplitudes [1958] = 8'd123;
   assign soundFileAmplitudes [1959] = 8'd130;
   assign soundFileAmplitudes [1960] = 8'd129;
   assign soundFileAmplitudes [1961] = 8'd121;
   assign soundFileAmplitudes [1962] = 8'd116;
   assign soundFileAmplitudes [1963] = 8'd108;
   assign soundFileAmplitudes [1964] = 8'd115;
   assign soundFileAmplitudes [1965] = 8'd120;
   assign soundFileAmplitudes [1966] = 8'd124;
   assign soundFileAmplitudes [1967] = 8'd140;
   assign soundFileAmplitudes [1968] = 8'd148;
   assign soundFileAmplitudes [1969] = 8'd140;
   assign soundFileAmplitudes [1970] = 8'd133;
   assign soundFileAmplitudes [1971] = 8'd127;
   assign soundFileAmplitudes [1972] = 8'd132;
   assign soundFileAmplitudes [1973] = 8'd134;
   assign soundFileAmplitudes [1974] = 8'd133;
   assign soundFileAmplitudes [1975] = 8'd137;
   assign soundFileAmplitudes [1976] = 8'd127;
   assign soundFileAmplitudes [1977] = 8'd124;
   assign soundFileAmplitudes [1978] = 8'd128;
   assign soundFileAmplitudes [1979] = 8'd135;
   assign soundFileAmplitudes [1980] = 8'd134;
   assign soundFileAmplitudes [1981] = 8'd132;
   assign soundFileAmplitudes [1982] = 8'd126;
   assign soundFileAmplitudes [1983] = 8'd123;
   assign soundFileAmplitudes [1984] = 8'd129;
   assign soundFileAmplitudes [1985] = 8'd117;
   assign soundFileAmplitudes [1986] = 8'd113;
   assign soundFileAmplitudes [1987] = 8'd113;
   assign soundFileAmplitudes [1988] = 8'd111;
   assign soundFileAmplitudes [1989] = 8'd113;
   assign soundFileAmplitudes [1990] = 8'd119;
   assign soundFileAmplitudes [1991] = 8'd125;
   assign soundFileAmplitudes [1992] = 8'd121;
   assign soundFileAmplitudes [1993] = 8'd118;
   assign soundFileAmplitudes [1994] = 8'd110;
   assign soundFileAmplitudes [1995] = 8'd120;
   assign soundFileAmplitudes [1996] = 8'd133;
   assign soundFileAmplitudes [1997] = 8'd133;
   assign soundFileAmplitudes [1998] = 8'd138;
   assign soundFileAmplitudes [1999] = 8'd139;
   assign soundFileAmplitudes [2000] = 8'd149;
   assign soundFileAmplitudes [2001] = 8'd139;
   assign soundFileAmplitudes [2002] = 8'd131;
   assign soundFileAmplitudes [2003] = 8'd136;
   assign soundFileAmplitudes [2004] = 8'd132;
   assign soundFileAmplitudes [2005] = 8'd133;
   assign soundFileAmplitudes [2006] = 8'd124;
   assign soundFileAmplitudes [2007] = 8'd117;
   assign soundFileAmplitudes [2008] = 8'd109;
   assign soundFileAmplitudes [2009] = 8'd100;
   assign soundFileAmplitudes [2010] = 8'd103;
   assign soundFileAmplitudes [2011] = 8'd109;
   assign soundFileAmplitudes [2012] = 8'd118;
   assign soundFileAmplitudes [2013] = 8'd133;
   assign soundFileAmplitudes [2014] = 8'd141;
   assign soundFileAmplitudes [2015] = 8'd144;
   assign soundFileAmplitudes [2016] = 8'd147;
   assign soundFileAmplitudes [2017] = 8'd146;
   assign soundFileAmplitudes [2018] = 8'd141;
   assign soundFileAmplitudes [2019] = 8'd138;
   assign soundFileAmplitudes [2020] = 8'd138;
   assign soundFileAmplitudes [2021] = 8'd136;
   assign soundFileAmplitudes [2022] = 8'd137;
   assign soundFileAmplitudes [2023] = 8'd129;
   assign soundFileAmplitudes [2024] = 8'd118;
   assign soundFileAmplitudes [2025] = 8'd112;
   assign soundFileAmplitudes [2026] = 8'd108;
   assign soundFileAmplitudes [2027] = 8'd106;
   assign soundFileAmplitudes [2028] = 8'd101;
   assign soundFileAmplitudes [2029] = 8'd102;
   assign soundFileAmplitudes [2030] = 8'd106;
   assign soundFileAmplitudes [2031] = 8'd117;
   assign soundFileAmplitudes [2032] = 8'd129;
   assign soundFileAmplitudes [2033] = 8'd136;
   assign soundFileAmplitudes [2034] = 8'd147;
   assign soundFileAmplitudes [2035] = 8'd149;
   assign soundFileAmplitudes [2036] = 8'd145;
   assign soundFileAmplitudes [2037] = 8'd135;
   assign soundFileAmplitudes [2038] = 8'd133;
   assign soundFileAmplitudes [2039] = 8'd126;
   assign soundFileAmplitudes [2040] = 8'd110;
   assign soundFileAmplitudes [2041] = 8'd104;
   assign soundFileAmplitudes [2042] = 8'd103;
   assign soundFileAmplitudes [2043] = 8'd114;
   assign soundFileAmplitudes [2044] = 8'd115;
   assign soundFileAmplitudes [2045] = 8'd112;
   assign soundFileAmplitudes [2046] = 8'd110;
   assign soundFileAmplitudes [2047] = 8'd111;
   assign soundFileAmplitudes [2048] = 8'd120;
   assign soundFileAmplitudes [2049] = 8'd133;
   assign soundFileAmplitudes [2050] = 8'd148;
   assign soundFileAmplitudes [2051] = 8'd151;
   assign soundFileAmplitudes [2052] = 8'd154;
   assign soundFileAmplitudes [2053] = 8'd155;
   assign soundFileAmplitudes [2054] = 8'd148;
   assign soundFileAmplitudes [2055] = 8'd145;
   assign soundFileAmplitudes [2056] = 8'd142;
   assign soundFileAmplitudes [2057] = 8'd140;
   assign soundFileAmplitudes [2058] = 8'd135;
   assign soundFileAmplitudes [2059] = 8'd127;
   assign soundFileAmplitudes [2060] = 8'd120;
   assign soundFileAmplitudes [2061] = 8'd104;
   assign soundFileAmplitudes [2062] = 8'd98;
   assign soundFileAmplitudes [2063] = 8'd101;
   assign soundFileAmplitudes [2064] = 8'd107;
   assign soundFileAmplitudes [2065] = 8'd114;
   assign soundFileAmplitudes [2066] = 8'd118;
   assign soundFileAmplitudes [2067] = 8'd125;
   assign soundFileAmplitudes [2068] = 8'd130;
   assign soundFileAmplitudes [2069] = 8'd127;
   assign soundFileAmplitudes [2070] = 8'd135;
   assign soundFileAmplitudes [2071] = 8'd138;
   assign soundFileAmplitudes [2072] = 8'd137;
   assign soundFileAmplitudes [2073] = 8'd130;
   assign soundFileAmplitudes [2074] = 8'd124;
   assign soundFileAmplitudes [2075] = 8'd125;
   assign soundFileAmplitudes [2076] = 8'd116;
   assign soundFileAmplitudes [2077] = 8'd115;
   assign soundFileAmplitudes [2078] = 8'd108;
   assign soundFileAmplitudes [2079] = 8'd109;
   assign soundFileAmplitudes [2080] = 8'd105;
   assign soundFileAmplitudes [2081] = 8'd105;
   assign soundFileAmplitudes [2082] = 8'd108;
   assign soundFileAmplitudes [2083] = 8'd116;
   assign soundFileAmplitudes [2084] = 8'd137;
   assign soundFileAmplitudes [2085] = 8'd149;
   assign soundFileAmplitudes [2086] = 8'd152;
   assign soundFileAmplitudes [2087] = 8'd151;
   assign soundFileAmplitudes [2088] = 8'd156;
   assign soundFileAmplitudes [2089] = 8'd155;
   assign soundFileAmplitudes [2090] = 8'd149;
   assign soundFileAmplitudes [2091] = 8'd149;
   assign soundFileAmplitudes [2092] = 8'd147;
   assign soundFileAmplitudes [2093] = 8'd143;
   assign soundFileAmplitudes [2094] = 8'd145;
   assign soundFileAmplitudes [2095] = 8'd139;
   assign soundFileAmplitudes [2096] = 8'd128;
   assign soundFileAmplitudes [2097] = 8'd119;
   assign soundFileAmplitudes [2098] = 8'd115;
   assign soundFileAmplitudes [2099] = 8'd113;
   assign soundFileAmplitudes [2100] = 8'd108;
   assign soundFileAmplitudes [2101] = 8'd97;
   assign soundFileAmplitudes [2102] = 8'd93;
   assign soundFileAmplitudes [2103] = 8'd93;
   assign soundFileAmplitudes [2104] = 8'd99;
   assign soundFileAmplitudes [2105] = 8'd108;
   assign soundFileAmplitudes [2106] = 8'd119;
   assign soundFileAmplitudes [2107] = 8'd130;
   assign soundFileAmplitudes [2108] = 8'd121;
   assign soundFileAmplitudes [2109] = 8'd115;
   assign soundFileAmplitudes [2110] = 8'd118;
   assign soundFileAmplitudes [2111] = 8'd115;
   assign soundFileAmplitudes [2112] = 8'd127;
   assign soundFileAmplitudes [2113] = 8'd130;
   assign soundFileAmplitudes [2114] = 8'd125;
   assign soundFileAmplitudes [2115] = 8'd125;
   assign soundFileAmplitudes [2116] = 8'd117;
   assign soundFileAmplitudes [2117] = 8'd103;
   assign soundFileAmplitudes [2118] = 8'd79;
   assign soundFileAmplitudes [2119] = 8'd107;
   assign soundFileAmplitudes [2120] = 8'd150;
   assign soundFileAmplitudes [2121] = 8'd149;
   assign soundFileAmplitudes [2122] = 8'd155;
   assign soundFileAmplitudes [2123] = 8'd164;
   assign soundFileAmplitudes [2124] = 8'd151;
   assign soundFileAmplitudes [2125] = 8'd155;
   assign soundFileAmplitudes [2126] = 8'd159;
   assign soundFileAmplitudes [2127] = 8'd160;
   assign soundFileAmplitudes [2128] = 8'd166;
   assign soundFileAmplitudes [2129] = 8'd155;
   assign soundFileAmplitudes [2130] = 8'd148;
   assign soundFileAmplitudes [2131] = 8'd140;
   assign soundFileAmplitudes [2132] = 8'd132;
   assign soundFileAmplitudes [2133] = 8'd121;
   assign soundFileAmplitudes [2134] = 8'd110;
   assign soundFileAmplitudes [2135] = 8'd96;
   assign soundFileAmplitudes [2136] = 8'd87;
   assign soundFileAmplitudes [2137] = 8'd83;
   assign soundFileAmplitudes [2138] = 8'd88;
   assign soundFileAmplitudes [2139] = 8'd92;
   assign soundFileAmplitudes [2140] = 8'd100;
   assign soundFileAmplitudes [2141] = 8'd111;
   assign soundFileAmplitudes [2142] = 8'd121;
   assign soundFileAmplitudes [2143] = 8'd112;
   assign soundFileAmplitudes [2144] = 8'd118;
   assign soundFileAmplitudes [2145] = 8'd133;
   assign soundFileAmplitudes [2146] = 8'd132;
   assign soundFileAmplitudes [2147] = 8'd138;
   assign soundFileAmplitudes [2148] = 8'd125;
   assign soundFileAmplitudes [2149] = 8'd121;
   assign soundFileAmplitudes [2150] = 8'd124;
   assign soundFileAmplitudes [2151] = 8'd124;
   assign soundFileAmplitudes [2152] = 8'd91;
   assign soundFileAmplitudes [2153] = 8'd121;
   assign soundFileAmplitudes [2154] = 8'd159;
   assign soundFileAmplitudes [2155] = 8'd148;
   assign soundFileAmplitudes [2156] = 8'd161;
   assign soundFileAmplitudes [2157] = 8'd163;
   assign soundFileAmplitudes [2158] = 8'd156;
   assign soundFileAmplitudes [2159] = 8'd165;
   assign soundFileAmplitudes [2160] = 8'd166;
   assign soundFileAmplitudes [2161] = 8'd148;
   assign soundFileAmplitudes [2162] = 8'd141;
   assign soundFileAmplitudes [2163] = 8'd132;
   assign soundFileAmplitudes [2164] = 8'd135;
   assign soundFileAmplitudes [2165] = 8'd128;
   assign soundFileAmplitudes [2166] = 8'd113;
   assign soundFileAmplitudes [2167] = 8'd92;
   assign soundFileAmplitudes [2168] = 8'd89;
   assign soundFileAmplitudes [2169] = 8'd97;
   assign soundFileAmplitudes [2170] = 8'd99;
   assign soundFileAmplitudes [2171] = 8'd103;
   assign soundFileAmplitudes [2172] = 8'd104;
   assign soundFileAmplitudes [2173] = 8'd96;
   assign soundFileAmplitudes [2174] = 8'd103;
   assign soundFileAmplitudes [2175] = 8'd117;
   assign soundFileAmplitudes [2176] = 8'd127;
   assign soundFileAmplitudes [2177] = 8'd130;
   assign soundFileAmplitudes [2178] = 8'd120;
   assign soundFileAmplitudes [2179] = 8'd125;
   assign soundFileAmplitudes [2180] = 8'd120;
   assign soundFileAmplitudes [2181] = 8'd105;
   assign soundFileAmplitudes [2182] = 8'd110;
   assign soundFileAmplitudes [2183] = 8'd115;
   assign soundFileAmplitudes [2184] = 8'd116;
   assign soundFileAmplitudes [2185] = 8'd117;
   assign soundFileAmplitudes [2186] = 8'd90;
   assign soundFileAmplitudes [2187] = 8'd118;
   assign soundFileAmplitudes [2188] = 8'd160;
   assign soundFileAmplitudes [2189] = 8'd168;
   assign soundFileAmplitudes [2190] = 8'd184;
   assign soundFileAmplitudes [2191] = 8'd193;
   assign soundFileAmplitudes [2192] = 8'd184;
   assign soundFileAmplitudes [2193] = 8'd177;
   assign soundFileAmplitudes [2194] = 8'd169;
   assign soundFileAmplitudes [2195] = 8'd161;
   assign soundFileAmplitudes [2196] = 8'd150;
   assign soundFileAmplitudes [2197] = 8'd129;
   assign soundFileAmplitudes [2198] = 8'd117;
   assign soundFileAmplitudes [2199] = 8'd107;
   assign soundFileAmplitudes [2200] = 8'd96;
   assign soundFileAmplitudes [2201] = 8'd83;
   assign soundFileAmplitudes [2202] = 8'd79;
   assign soundFileAmplitudes [2203] = 8'd85;
   assign soundFileAmplitudes [2204] = 8'd85;
   assign soundFileAmplitudes [2205] = 8'd92;
   assign soundFileAmplitudes [2206] = 8'd107;
   assign soundFileAmplitudes [2207] = 8'd110;
   assign soundFileAmplitudes [2208] = 8'd116;
   assign soundFileAmplitudes [2209] = 8'd130;
   assign soundFileAmplitudes [2210] = 8'd143;
   assign soundFileAmplitudes [2211] = 8'd142;
   assign soundFileAmplitudes [2212] = 8'd144;
   assign soundFileAmplitudes [2213] = 8'd123;
   assign soundFileAmplitudes [2214] = 8'd109;
   assign soundFileAmplitudes [2215] = 8'd116;
   assign soundFileAmplitudes [2216] = 8'd119;
   assign soundFileAmplitudes [2217] = 8'd121;
   assign soundFileAmplitudes [2218] = 8'd113;
   assign soundFileAmplitudes [2219] = 8'd106;
   assign soundFileAmplitudes [2220] = 8'd96;
   assign soundFileAmplitudes [2221] = 8'd113;
   assign soundFileAmplitudes [2222] = 8'd139;
   assign soundFileAmplitudes [2223] = 8'd162;
   assign soundFileAmplitudes [2224] = 8'd176;
   assign soundFileAmplitudes [2225] = 8'd181;
   assign soundFileAmplitudes [2226] = 8'd182;
   assign soundFileAmplitudes [2227] = 8'd173;
   assign soundFileAmplitudes [2228] = 8'd165;
   assign soundFileAmplitudes [2229] = 8'd160;
   assign soundFileAmplitudes [2230] = 8'd153;
   assign soundFileAmplitudes [2231] = 8'd132;
   assign soundFileAmplitudes [2232] = 8'd114;
   assign soundFileAmplitudes [2233] = 8'd117;
   assign soundFileAmplitudes [2234] = 8'd109;
   assign soundFileAmplitudes [2235] = 8'd92;
   assign soundFileAmplitudes [2236] = 8'd78;
   assign soundFileAmplitudes [2237] = 8'd69;
   assign soundFileAmplitudes [2238] = 8'd86;
   assign soundFileAmplitudes [2239] = 8'd90;
   assign soundFileAmplitudes [2240] = 8'd92;
   assign soundFileAmplitudes [2241] = 8'd98;
   assign soundFileAmplitudes [2242] = 8'd109;
   assign soundFileAmplitudes [2243] = 8'd124;
   assign soundFileAmplitudes [2244] = 8'd125;
   assign soundFileAmplitudes [2245] = 8'd131;
   assign soundFileAmplitudes [2246] = 8'd136;
   assign soundFileAmplitudes [2247] = 8'd139;
   assign soundFileAmplitudes [2248] = 8'd126;
   assign soundFileAmplitudes [2249] = 8'd120;
   assign soundFileAmplitudes [2250] = 8'd115;
   assign soundFileAmplitudes [2251] = 8'd115;
   assign soundFileAmplitudes [2252] = 8'd134;
   assign soundFileAmplitudes [2253] = 8'd149;
   assign soundFileAmplitudes [2254] = 8'd145;
   assign soundFileAmplitudes [2255] = 8'd125;
   assign soundFileAmplitudes [2256] = 8'd123;
   assign soundFileAmplitudes [2257] = 8'd140;
   assign soundFileAmplitudes [2258] = 8'd155;
   assign soundFileAmplitudes [2259] = 8'd153;
   assign soundFileAmplitudes [2260] = 8'd152;
   assign soundFileAmplitudes [2261] = 8'd150;
   assign soundFileAmplitudes [2262] = 8'd145;
   assign soundFileAmplitudes [2263] = 8'd152;
   assign soundFileAmplitudes [2264] = 8'd155;
   assign soundFileAmplitudes [2265] = 8'd150;
   assign soundFileAmplitudes [2266] = 8'd146;
   assign soundFileAmplitudes [2267] = 8'd132;
   assign soundFileAmplitudes [2268] = 8'd123;
   assign soundFileAmplitudes [2269] = 8'd122;
   assign soundFileAmplitudes [2270] = 8'd115;
   assign soundFileAmplitudes [2271] = 8'd106;
   assign soundFileAmplitudes [2272] = 8'd106;
   assign soundFileAmplitudes [2273] = 8'd97;
   assign soundFileAmplitudes [2274] = 8'd103;
   assign soundFileAmplitudes [2275] = 8'd100;
   assign soundFileAmplitudes [2276] = 8'd87;
   assign soundFileAmplitudes [2277] = 8'd94;
   assign soundFileAmplitudes [2278] = 8'd103;
   assign soundFileAmplitudes [2279] = 8'd110;
   assign soundFileAmplitudes [2280] = 8'd111;
   assign soundFileAmplitudes [2281] = 8'd119;
   assign soundFileAmplitudes [2282] = 8'd130;
   assign soundFileAmplitudes [2283] = 8'd123;
   assign soundFileAmplitudes [2284] = 8'd119;
   assign soundFileAmplitudes [2285] = 8'd131;
   assign soundFileAmplitudes [2286] = 8'd126;
   assign soundFileAmplitudes [2287] = 8'd133;
   assign soundFileAmplitudes [2288] = 8'd131;
   assign soundFileAmplitudes [2289] = 8'd122;
   assign soundFileAmplitudes [2290] = 8'd125;
   assign soundFileAmplitudes [2291] = 8'd128;
   assign soundFileAmplitudes [2292] = 8'd133;
   assign soundFileAmplitudes [2293] = 8'd136;
   assign soundFileAmplitudes [2294] = 8'd135;
   assign soundFileAmplitudes [2295] = 8'd137;
   assign soundFileAmplitudes [2296] = 8'd146;
   assign soundFileAmplitudes [2297] = 8'd155;
   assign soundFileAmplitudes [2298] = 8'd158;
   assign soundFileAmplitudes [2299] = 8'd153;
   assign soundFileAmplitudes [2300] = 8'd148;
   assign soundFileAmplitudes [2301] = 8'd142;
   assign soundFileAmplitudes [2302] = 8'd137;
   assign soundFileAmplitudes [2303] = 8'd133;
   assign soundFileAmplitudes [2304] = 8'd123;
   assign soundFileAmplitudes [2305] = 8'd125;
   assign soundFileAmplitudes [2306] = 8'd118;
   assign soundFileAmplitudes [2307] = 8'd107;
   assign soundFileAmplitudes [2308] = 8'd110;
   assign soundFileAmplitudes [2309] = 8'd108;
   assign soundFileAmplitudes [2310] = 8'd114;
   assign soundFileAmplitudes [2311] = 8'd115;
   assign soundFileAmplitudes [2312] = 8'd110;
   assign soundFileAmplitudes [2313] = 8'd108;
   assign soundFileAmplitudes [2314] = 8'd109;
   assign soundFileAmplitudes [2315] = 8'd110;
   assign soundFileAmplitudes [2316] = 8'd124;
   assign soundFileAmplitudes [2317] = 8'd137;
   assign soundFileAmplitudes [2318] = 8'd127;
   assign soundFileAmplitudes [2319] = 8'd114;
   assign soundFileAmplitudes [2320] = 8'd106;
   assign soundFileAmplitudes [2321] = 8'd101;
   assign soundFileAmplitudes [2322] = 8'd99;
   assign soundFileAmplitudes [2323] = 8'd105;
   assign soundFileAmplitudes [2324] = 8'd107;
   assign soundFileAmplitudes [2325] = 8'd110;
   assign soundFileAmplitudes [2326] = 8'd116;
   assign soundFileAmplitudes [2327] = 8'd123;
   assign soundFileAmplitudes [2328] = 8'd140;
   assign soundFileAmplitudes [2329] = 8'd155;
   assign soundFileAmplitudes [2330] = 8'd166;
   assign soundFileAmplitudes [2331] = 8'd177;
   assign soundFileAmplitudes [2332] = 8'd174;
   assign soundFileAmplitudes [2333] = 8'd173;
   assign soundFileAmplitudes [2334] = 8'd177;
   assign soundFileAmplitudes [2335] = 8'd169;
   assign soundFileAmplitudes [2336] = 8'd155;
   assign soundFileAmplitudes [2337] = 8'd145;
   assign soundFileAmplitudes [2338] = 8'd131;
   assign soundFileAmplitudes [2339] = 8'd113;
   assign soundFileAmplitudes [2340] = 8'd109;
   assign soundFileAmplitudes [2341] = 8'd103;
   assign soundFileAmplitudes [2342] = 8'd105;
   assign soundFileAmplitudes [2343] = 8'd105;
   assign soundFileAmplitudes [2344] = 8'd102;
   assign soundFileAmplitudes [2345] = 8'd99;
   assign soundFileAmplitudes [2346] = 8'd91;
   assign soundFileAmplitudes [2347] = 8'd100;
   assign soundFileAmplitudes [2348] = 8'd118;
   assign soundFileAmplitudes [2349] = 8'd138;
   assign soundFileAmplitudes [2350] = 8'd132;
   assign soundFileAmplitudes [2351] = 8'd121;
   assign soundFileAmplitudes [2352] = 8'd116;
   assign soundFileAmplitudes [2353] = 8'd105;
   assign soundFileAmplitudes [2354] = 8'd95;
   assign soundFileAmplitudes [2355] = 8'd90;
   assign soundFileAmplitudes [2356] = 8'd98;
   assign soundFileAmplitudes [2357] = 8'd101;
   assign soundFileAmplitudes [2358] = 8'd97;
   assign soundFileAmplitudes [2359] = 8'd97;
   assign soundFileAmplitudes [2360] = 8'd101;
   assign soundFileAmplitudes [2361] = 8'd123;
   assign soundFileAmplitudes [2362] = 8'd144;
   assign soundFileAmplitudes [2363] = 8'd165;
   assign soundFileAmplitudes [2364] = 8'd179;
   assign soundFileAmplitudes [2365] = 8'd172;
   assign soundFileAmplitudes [2366] = 8'd177;
   assign soundFileAmplitudes [2367] = 8'd186;
   assign soundFileAmplitudes [2368] = 8'd184;
   assign soundFileAmplitudes [2369] = 8'd180;
   assign soundFileAmplitudes [2370] = 8'd175;
   assign soundFileAmplitudes [2371] = 8'd154;
   assign soundFileAmplitudes [2372] = 8'd133;
   assign soundFileAmplitudes [2373] = 8'd123;
   assign soundFileAmplitudes [2374] = 8'd112;
   assign soundFileAmplitudes [2375] = 8'd103;
   assign soundFileAmplitudes [2376] = 8'd99;
   assign soundFileAmplitudes [2377] = 8'd92;
   assign soundFileAmplitudes [2378] = 8'd88;
   assign soundFileAmplitudes [2379] = 8'd92;
   assign soundFileAmplitudes [2380] = 8'd95;
   assign soundFileAmplitudes [2381] = 8'd109;
   assign soundFileAmplitudes [2382] = 8'd106;
   assign soundFileAmplitudes [2383] = 8'd102;
   assign soundFileAmplitudes [2384] = 8'd105;
   assign soundFileAmplitudes [2385] = 8'd117;
   assign soundFileAmplitudes [2386] = 8'd127;
   assign soundFileAmplitudes [2387] = 8'd113;
   assign soundFileAmplitudes [2388] = 8'd110;
   assign soundFileAmplitudes [2389] = 8'd95;
   assign soundFileAmplitudes [2390] = 8'd94;
   assign soundFileAmplitudes [2391] = 8'd102;
   assign soundFileAmplitudes [2392] = 8'd94;
   assign soundFileAmplitudes [2393] = 8'd102;
   assign soundFileAmplitudes [2394] = 8'd113;
   assign soundFileAmplitudes [2395] = 8'd118;
   assign soundFileAmplitudes [2396] = 8'd140;
   assign soundFileAmplitudes [2397] = 8'd157;
   assign soundFileAmplitudes [2398] = 8'd158;
   assign soundFileAmplitudes [2399] = 8'd164;
   assign soundFileAmplitudes [2400] = 8'd169;
   assign soundFileAmplitudes [2401] = 8'd185;
   assign soundFileAmplitudes [2402] = 8'd199;
   assign soundFileAmplitudes [2403] = 8'd191;
   assign soundFileAmplitudes [2404] = 8'd175;
   assign soundFileAmplitudes [2405] = 8'd163;
   assign soundFileAmplitudes [2406] = 8'd147;
   assign soundFileAmplitudes [2407] = 8'd136;
   assign soundFileAmplitudes [2408] = 8'd128;
   assign soundFileAmplitudes [2409] = 8'd116;
   assign soundFileAmplitudes [2410] = 8'd112;
   assign soundFileAmplitudes [2411] = 8'd109;
   assign soundFileAmplitudes [2412] = 8'd105;
   assign soundFileAmplitudes [2413] = 8'd105;
   assign soundFileAmplitudes [2414] = 8'd104;
   assign soundFileAmplitudes [2415] = 8'd95;
   assign soundFileAmplitudes [2416] = 8'd87;
   assign soundFileAmplitudes [2417] = 8'd83;
   assign soundFileAmplitudes [2418] = 8'd91;
   assign soundFileAmplitudes [2419] = 8'd105;
   assign soundFileAmplitudes [2420] = 8'd119;
   assign soundFileAmplitudes [2421] = 8'd118;
   assign soundFileAmplitudes [2422] = 8'd112;
   assign soundFileAmplitudes [2423] = 8'd115;
   assign soundFileAmplitudes [2424] = 8'd119;
   assign soundFileAmplitudes [2425] = 8'd117;
   assign soundFileAmplitudes [2426] = 8'd114;
   assign soundFileAmplitudes [2427] = 8'd119;
   assign soundFileAmplitudes [2428] = 8'd111;
   assign soundFileAmplitudes [2429] = 8'd122;
   assign soundFileAmplitudes [2430] = 8'd135;
   assign soundFileAmplitudes [2431] = 8'd137;
   assign soundFileAmplitudes [2432] = 8'd145;
   assign soundFileAmplitudes [2433] = 8'd157;
   assign soundFileAmplitudes [2434] = 8'd163;
   assign soundFileAmplitudes [2435] = 8'd157;
   assign soundFileAmplitudes [2436] = 8'd151;
   assign soundFileAmplitudes [2437] = 8'd149;
   assign soundFileAmplitudes [2438] = 8'd151;
   assign soundFileAmplitudes [2439] = 8'd150;
   assign soundFileAmplitudes [2440] = 8'd139;
   assign soundFileAmplitudes [2441] = 8'd140;
   assign soundFileAmplitudes [2442] = 8'd133;
   assign soundFileAmplitudes [2443] = 8'd125;
   assign soundFileAmplitudes [2444] = 8'd117;
   assign soundFileAmplitudes [2445] = 8'd117;
   assign soundFileAmplitudes [2446] = 8'd135;
   assign soundFileAmplitudes [2447] = 8'd123;
   assign soundFileAmplitudes [2448] = 8'd114;
   assign soundFileAmplitudes [2449] = 8'd102;
   assign soundFileAmplitudes [2450] = 8'd98;
   assign soundFileAmplitudes [2451] = 8'd101;
   assign soundFileAmplitudes [2452] = 8'd103;
   assign soundFileAmplitudes [2453] = 8'd99;
   assign soundFileAmplitudes [2454] = 8'd93;
   assign soundFileAmplitudes [2455] = 8'd94;
   assign soundFileAmplitudes [2456] = 8'd108;
   assign soundFileAmplitudes [2457] = 8'd121;
   assign soundFileAmplitudes [2458] = 8'd133;
   assign soundFileAmplitudes [2459] = 8'd147;
   assign soundFileAmplitudes [2460] = 8'd141;
   assign soundFileAmplitudes [2461] = 8'd143;
   assign soundFileAmplitudes [2462] = 8'd138;
   assign soundFileAmplitudes [2463] = 8'd139;
   assign soundFileAmplitudes [2464] = 8'd139;
   assign soundFileAmplitudes [2465] = 8'd140;
   assign soundFileAmplitudes [2466] = 8'd137;
   assign soundFileAmplitudes [2467] = 8'd142;
   assign soundFileAmplitudes [2468] = 8'd141;
   assign soundFileAmplitudes [2469] = 8'd126;
   assign soundFileAmplitudes [2470] = 8'd119;
   assign soundFileAmplitudes [2471] = 8'd108;
   assign soundFileAmplitudes [2472] = 8'd111;
   assign soundFileAmplitudes [2473] = 8'd130;
   assign soundFileAmplitudes [2474] = 8'd140;
   assign soundFileAmplitudes [2475] = 8'd137;
   assign soundFileAmplitudes [2476] = 8'd138;
   assign soundFileAmplitudes [2477] = 8'd129;
   assign soundFileAmplitudes [2478] = 8'd131;
   assign soundFileAmplitudes [2479] = 8'd137;
   assign soundFileAmplitudes [2480] = 8'd134;
   assign soundFileAmplitudes [2481] = 8'd136;
   assign soundFileAmplitudes [2482] = 8'd130;
   assign soundFileAmplitudes [2483] = 8'd121;
   assign soundFileAmplitudes [2484] = 8'd119;
   assign soundFileAmplitudes [2485] = 8'd118;
   assign soundFileAmplitudes [2486] = 8'd112;
   assign soundFileAmplitudes [2487] = 8'd96;
   assign soundFileAmplitudes [2488] = 8'd88;
   assign soundFileAmplitudes [2489] = 8'd98;
   assign soundFileAmplitudes [2490] = 8'd111;
   assign soundFileAmplitudes [2491] = 8'd121;
   assign soundFileAmplitudes [2492] = 8'd127;
   assign soundFileAmplitudes [2493] = 8'd125;
   assign soundFileAmplitudes [2494] = 8'd134;
   assign soundFileAmplitudes [2495] = 8'd143;
   assign soundFileAmplitudes [2496] = 8'd138;
   assign soundFileAmplitudes [2497] = 8'd144;
   assign soundFileAmplitudes [2498] = 8'd141;
   assign soundFileAmplitudes [2499] = 8'd132;
   assign soundFileAmplitudes [2500] = 8'd124;
   assign soundFileAmplitudes [2501] = 8'd122;
   assign soundFileAmplitudes [2502] = 8'd121;
   assign soundFileAmplitudes [2503] = 8'd124;
   assign soundFileAmplitudes [2504] = 8'd122;
   assign soundFileAmplitudes [2505] = 8'd114;
   assign soundFileAmplitudes [2506] = 8'd109;
   assign soundFileAmplitudes [2507] = 8'd118;
   assign soundFileAmplitudes [2508] = 8'd122;
   assign soundFileAmplitudes [2509] = 8'd125;
   assign soundFileAmplitudes [2510] = 8'd130;
   assign soundFileAmplitudes [2511] = 8'd130;
   assign soundFileAmplitudes [2512] = 8'd143;
   assign soundFileAmplitudes [2513] = 8'd139;
   assign soundFileAmplitudes [2514] = 8'd132;
   assign soundFileAmplitudes [2515] = 8'd125;
   assign soundFileAmplitudes [2516] = 8'd124;
   assign soundFileAmplitudes [2517] = 8'd132;
   assign soundFileAmplitudes [2518] = 8'd133;
   assign soundFileAmplitudes [2519] = 8'd131;
   assign soundFileAmplitudes [2520] = 8'd125;
   assign soundFileAmplitudes [2521] = 8'd121;
   assign soundFileAmplitudes [2522] = 8'd120;
   assign soundFileAmplitudes [2523] = 8'd117;
   assign soundFileAmplitudes [2524] = 8'd113;
   assign soundFileAmplitudes [2525] = 8'd109;
   assign soundFileAmplitudes [2526] = 8'd109;
   assign soundFileAmplitudes [2527] = 8'd122;
   assign soundFileAmplitudes [2528] = 8'd134;
   assign soundFileAmplitudes [2529] = 8'd153;
   assign soundFileAmplitudes [2530] = 8'd159;
   assign soundFileAmplitudes [2531] = 8'd143;
   assign soundFileAmplitudes [2532] = 8'd126;
   assign soundFileAmplitudes [2533] = 8'd121;
   assign soundFileAmplitudes [2534] = 8'd116;
   assign soundFileAmplitudes [2535] = 8'd118;
   assign soundFileAmplitudes [2536] = 8'd120;
   assign soundFileAmplitudes [2537] = 8'd112;
   assign soundFileAmplitudes [2538] = 8'd114;
   assign soundFileAmplitudes [2539] = 8'd112;
   assign soundFileAmplitudes [2540] = 8'd114;
   assign soundFileAmplitudes [2541] = 8'd128;
   assign soundFileAmplitudes [2542] = 8'd130;
   assign soundFileAmplitudes [2543] = 8'd130;
   assign soundFileAmplitudes [2544] = 8'd141;
   assign soundFileAmplitudes [2545] = 8'd150;
   assign soundFileAmplitudes [2546] = 8'd145;
   assign soundFileAmplitudes [2547] = 8'd137;
   assign soundFileAmplitudes [2548] = 8'd123;
   assign soundFileAmplitudes [2549] = 8'd123;
   assign soundFileAmplitudes [2550] = 8'd126;
   assign soundFileAmplitudes [2551] = 8'd130;
   assign soundFileAmplitudes [2552] = 8'd139;
   assign soundFileAmplitudes [2553] = 8'd137;
   assign soundFileAmplitudes [2554] = 8'd129;
   assign soundFileAmplitudes [2555] = 8'd122;
   assign soundFileAmplitudes [2556] = 8'd123;
   assign soundFileAmplitudes [2557] = 8'd118;
   assign soundFileAmplitudes [2558] = 8'd108;
   assign soundFileAmplitudes [2559] = 8'd107;
   assign soundFileAmplitudes [2560] = 8'd121;
   assign soundFileAmplitudes [2561] = 8'd125;
   assign soundFileAmplitudes [2562] = 8'd128;
   assign soundFileAmplitudes [2563] = 8'd137;
   assign soundFileAmplitudes [2564] = 8'd139;
   assign soundFileAmplitudes [2565] = 8'd141;
   assign soundFileAmplitudes [2566] = 8'd140;
   assign soundFileAmplitudes [2567] = 8'd130;
   assign soundFileAmplitudes [2568] = 8'd111;
   assign soundFileAmplitudes [2569] = 8'd93;
   assign soundFileAmplitudes [2570] = 8'd87;
   assign soundFileAmplitudes [2571] = 8'd89;
   assign soundFileAmplitudes [2572] = 8'd94;
   assign soundFileAmplitudes [2573] = 8'd105;
   assign soundFileAmplitudes [2574] = 8'd112;
   assign soundFileAmplitudes [2575] = 8'd119;
   assign soundFileAmplitudes [2576] = 8'd136;
   assign soundFileAmplitudes [2577] = 8'd148;
   assign soundFileAmplitudes [2578] = 8'd149;
   assign soundFileAmplitudes [2579] = 8'd151;
   assign soundFileAmplitudes [2580] = 8'd153;
   assign soundFileAmplitudes [2581] = 8'd155;
   assign soundFileAmplitudes [2582] = 8'd160;
   assign soundFileAmplitudes [2583] = 8'd154;
   assign soundFileAmplitudes [2584] = 8'd136;
   assign soundFileAmplitudes [2585] = 8'd121;
   assign soundFileAmplitudes [2586] = 8'd107;
   assign soundFileAmplitudes [2587] = 8'd108;
   assign soundFileAmplitudes [2588] = 8'd124;
   assign soundFileAmplitudes [2589] = 8'd132;
   assign soundFileAmplitudes [2590] = 8'd120;
   assign soundFileAmplitudes [2591] = 8'd118;
   assign soundFileAmplitudes [2592] = 8'd119;
   assign soundFileAmplitudes [2593] = 8'd121;
   assign soundFileAmplitudes [2594] = 8'd123;
   assign soundFileAmplitudes [2595] = 8'd128;
   assign soundFileAmplitudes [2596] = 8'd131;
   assign soundFileAmplitudes [2597] = 8'd133;
   assign soundFileAmplitudes [2598] = 8'd139;
   assign soundFileAmplitudes [2599] = 8'd137;
   assign soundFileAmplitudes [2600] = 8'd123;
   assign soundFileAmplitudes [2601] = 8'd115;
   assign soundFileAmplitudes [2602] = 8'd117;
   assign soundFileAmplitudes [2603] = 8'd106;
   assign soundFileAmplitudes [2604] = 8'd101;
   assign soundFileAmplitudes [2605] = 8'd101;
   assign soundFileAmplitudes [2606] = 8'd107;
   assign soundFileAmplitudes [2607] = 8'd110;
   assign soundFileAmplitudes [2608] = 8'd116;
   assign soundFileAmplitudes [2609] = 8'd120;
   assign soundFileAmplitudes [2610] = 8'd136;
   assign soundFileAmplitudes [2611] = 8'd146;
   assign soundFileAmplitudes [2612] = 8'd143;
   assign soundFileAmplitudes [2613] = 8'd147;
   assign soundFileAmplitudes [2614] = 8'd143;
   assign soundFileAmplitudes [2615] = 8'd143;
   assign soundFileAmplitudes [2616] = 8'd148;
   assign soundFileAmplitudes [2617] = 8'd150;
   assign soundFileAmplitudes [2618] = 8'd143;
   assign soundFileAmplitudes [2619] = 8'd143;
   assign soundFileAmplitudes [2620] = 8'd131;
   assign soundFileAmplitudes [2621] = 8'd122;
   assign soundFileAmplitudes [2622] = 8'd114;
   assign soundFileAmplitudes [2623] = 8'd111;
   assign soundFileAmplitudes [2624] = 8'd129;
   assign soundFileAmplitudes [2625] = 8'd130;
   assign soundFileAmplitudes [2626] = 8'd123;
   assign soundFileAmplitudes [2627] = 8'd118;
   assign soundFileAmplitudes [2628] = 8'd123;
   assign soundFileAmplitudes [2629] = 8'd129;
   assign soundFileAmplitudes [2630] = 8'd135;
   assign soundFileAmplitudes [2631] = 8'd131;
   assign soundFileAmplitudes [2632] = 8'd117;
   assign soundFileAmplitudes [2633] = 8'd102;
   assign soundFileAmplitudes [2634] = 8'd100;
   assign soundFileAmplitudes [2635] = 8'd112;
   assign soundFileAmplitudes [2636] = 8'd125;
   assign soundFileAmplitudes [2637] = 8'd126;
   assign soundFileAmplitudes [2638] = 8'd126;
   assign soundFileAmplitudes [2639] = 8'd118;
   assign soundFileAmplitudes [2640] = 8'd110;
   assign soundFileAmplitudes [2641] = 8'd109;
   assign soundFileAmplitudes [2642] = 8'd109;
   assign soundFileAmplitudes [2643] = 8'd122;
   assign soundFileAmplitudes [2644] = 8'd127;
   assign soundFileAmplitudes [2645] = 8'd125;
   assign soundFileAmplitudes [2646] = 8'd118;
   assign soundFileAmplitudes [2647] = 8'd117;
   assign soundFileAmplitudes [2648] = 8'd123;
   assign soundFileAmplitudes [2649] = 8'd131;
   assign soundFileAmplitudes [2650] = 8'd134;
   assign soundFileAmplitudes [2651] = 8'd141;
   assign soundFileAmplitudes [2652] = 8'd148;
   assign soundFileAmplitudes [2653] = 8'd146;
   assign soundFileAmplitudes [2654] = 8'd146;
   assign soundFileAmplitudes [2655] = 8'd148;
   assign soundFileAmplitudes [2656] = 8'd140;
   assign soundFileAmplitudes [2657] = 8'd142;
   assign soundFileAmplitudes [2658] = 8'd138;
   assign soundFileAmplitudes [2659] = 8'd124;
   assign soundFileAmplitudes [2660] = 8'd134;
   assign soundFileAmplitudes [2661] = 8'd135;
   assign soundFileAmplitudes [2662] = 8'd141;
   assign soundFileAmplitudes [2663] = 8'd132;
   assign soundFileAmplitudes [2664] = 8'd124;
   assign soundFileAmplitudes [2665] = 8'd112;
   assign soundFileAmplitudes [2666] = 8'd98;
   assign soundFileAmplitudes [2667] = 8'd107;
   assign soundFileAmplitudes [2668] = 8'd101;
   assign soundFileAmplitudes [2669] = 8'd98;
   assign soundFileAmplitudes [2670] = 8'd109;
   assign soundFileAmplitudes [2671] = 8'd105;
   assign soundFileAmplitudes [2672] = 8'd109;
   assign soundFileAmplitudes [2673] = 8'd120;
   assign soundFileAmplitudes [2674] = 8'd126;
   assign soundFileAmplitudes [2675] = 8'd124;
   assign soundFileAmplitudes [2676] = 8'd113;
   assign soundFileAmplitudes [2677] = 8'd117;
   assign soundFileAmplitudes [2678] = 8'd119;
   assign soundFileAmplitudes [2679] = 8'd128;
   assign soundFileAmplitudes [2680] = 8'd129;
   assign soundFileAmplitudes [2681] = 8'd128;
   assign soundFileAmplitudes [2682] = 8'd128;
   assign soundFileAmplitudes [2683] = 8'd132;
   assign soundFileAmplitudes [2684] = 8'd134;
   assign soundFileAmplitudes [2685] = 8'd132;
   assign soundFileAmplitudes [2686] = 8'd130;
   assign soundFileAmplitudes [2687] = 8'd132;
   assign soundFileAmplitudes [2688] = 8'd144;
   assign soundFileAmplitudes [2689] = 8'd150;
   assign soundFileAmplitudes [2690] = 8'd151;
   assign soundFileAmplitudes [2691] = 8'd142;
   assign soundFileAmplitudes [2692] = 8'd139;
   assign soundFileAmplitudes [2693] = 8'd140;
   assign soundFileAmplitudes [2694] = 8'd141;
   assign soundFileAmplitudes [2695] = 8'd141;
   assign soundFileAmplitudes [2696] = 8'd152;
   assign soundFileAmplitudes [2697] = 8'd142;
   assign soundFileAmplitudes [2698] = 8'd135;
   assign soundFileAmplitudes [2699] = 8'd118;
   assign soundFileAmplitudes [2700] = 8'd106;
   assign soundFileAmplitudes [2701] = 8'd110;
   assign soundFileAmplitudes [2702] = 8'd95;
   assign soundFileAmplitudes [2703] = 8'd97;
   assign soundFileAmplitudes [2704] = 8'd93;
   assign soundFileAmplitudes [2705] = 8'd95;
   assign soundFileAmplitudes [2706] = 8'd92;
   assign soundFileAmplitudes [2707] = 8'd96;
   assign soundFileAmplitudes [2708] = 8'd100;
   assign soundFileAmplitudes [2709] = 8'd110;
   assign soundFileAmplitudes [2710] = 8'd114;
   assign soundFileAmplitudes [2711] = 8'd112;
   assign soundFileAmplitudes [2712] = 8'd122;
   assign soundFileAmplitudes [2713] = 8'd130;
   assign soundFileAmplitudes [2714] = 8'd140;
   assign soundFileAmplitudes [2715] = 8'd144;
   assign soundFileAmplitudes [2716] = 8'd150;
   assign soundFileAmplitudes [2717] = 8'd143;
   assign soundFileAmplitudes [2718] = 8'd144;
   assign soundFileAmplitudes [2719] = 8'd153;
   assign soundFileAmplitudes [2720] = 8'd151;
   assign soundFileAmplitudes [2721] = 8'd147;
   assign soundFileAmplitudes [2722] = 8'd138;
   assign soundFileAmplitudes [2723] = 8'd129;
   assign soundFileAmplitudes [2724] = 8'd132;
   assign soundFileAmplitudes [2725] = 8'd145;
   assign soundFileAmplitudes [2726] = 8'd159;
   assign soundFileAmplitudes [2727] = 8'd168;
   assign soundFileAmplitudes [2728] = 8'd160;
   assign soundFileAmplitudes [2729] = 8'd153;
   assign soundFileAmplitudes [2730] = 8'd145;
   assign soundFileAmplitudes [2731] = 8'd117;
   assign soundFileAmplitudes [2732] = 8'd112;
   assign soundFileAmplitudes [2733] = 8'd116;
   assign soundFileAmplitudes [2734] = 8'd108;
   assign soundFileAmplitudes [2735] = 8'd102;
   assign soundFileAmplitudes [2736] = 8'd110;
   assign soundFileAmplitudes [2737] = 8'd107;
   assign soundFileAmplitudes [2738] = 8'd86;
   assign soundFileAmplitudes [2739] = 8'd82;
   assign soundFileAmplitudes [2740] = 8'd77;
   assign soundFileAmplitudes [2741] = 8'd84;
   assign soundFileAmplitudes [2742] = 8'd98;
   assign soundFileAmplitudes [2743] = 8'd102;
   assign soundFileAmplitudes [2744] = 8'd111;
   assign soundFileAmplitudes [2745] = 8'd114;
   assign soundFileAmplitudes [2746] = 8'd119;
   assign soundFileAmplitudes [2747] = 8'd126;
   assign soundFileAmplitudes [2748] = 8'd139;
   assign soundFileAmplitudes [2749] = 8'd140;
   assign soundFileAmplitudes [2750] = 8'd126;
   assign soundFileAmplitudes [2751] = 8'd133;
   assign soundFileAmplitudes [2752] = 8'd137;
   assign soundFileAmplitudes [2753] = 8'd138;
   assign soundFileAmplitudes [2754] = 8'd140;
   assign soundFileAmplitudes [2755] = 8'd154;
   assign soundFileAmplitudes [2756] = 8'd157;
   assign soundFileAmplitudes [2757] = 8'd157;
   assign soundFileAmplitudes [2758] = 8'd156;
   assign soundFileAmplitudes [2759] = 8'd142;
   assign soundFileAmplitudes [2760] = 8'd146;
   assign soundFileAmplitudes [2761] = 8'd163;
   assign soundFileAmplitudes [2762] = 8'd160;
   assign soundFileAmplitudes [2763] = 8'd153;
   assign soundFileAmplitudes [2764] = 8'd138;
   assign soundFileAmplitudes [2765] = 8'd121;
   assign soundFileAmplitudes [2766] = 8'd117;
   assign soundFileAmplitudes [2767] = 8'd92;
   assign soundFileAmplitudes [2768] = 8'd95;
   assign soundFileAmplitudes [2769] = 8'd116;
   assign soundFileAmplitudes [2770] = 8'd110;
   assign soundFileAmplitudes [2771] = 8'd109;
   assign soundFileAmplitudes [2772] = 8'd106;
   assign soundFileAmplitudes [2773] = 8'd104;
   assign soundFileAmplitudes [2774] = 8'd118;
   assign soundFileAmplitudes [2775] = 8'd119;
   assign soundFileAmplitudes [2776] = 8'd112;
   assign soundFileAmplitudes [2777] = 8'd110;
   assign soundFileAmplitudes [2778] = 8'd111;
   assign soundFileAmplitudes [2779] = 8'd111;
   assign soundFileAmplitudes [2780] = 8'd117;
   assign soundFileAmplitudes [2781] = 8'd119;
   assign soundFileAmplitudes [2782] = 8'd112;
   assign soundFileAmplitudes [2783] = 8'd109;
   assign soundFileAmplitudes [2784] = 8'd116;
   assign soundFileAmplitudes [2785] = 8'd125;
   assign soundFileAmplitudes [2786] = 8'd132;
   assign soundFileAmplitudes [2787] = 8'd138;
   assign soundFileAmplitudes [2788] = 8'd133;
   assign soundFileAmplitudes [2789] = 8'd133;
   assign soundFileAmplitudes [2790] = 8'd140;
   assign soundFileAmplitudes [2791] = 8'd139;
   assign soundFileAmplitudes [2792] = 8'd140;
   assign soundFileAmplitudes [2793] = 8'd147;
   assign soundFileAmplitudes [2794] = 8'd152;
   assign soundFileAmplitudes [2795] = 8'd152;
   assign soundFileAmplitudes [2796] = 8'd123;
   assign soundFileAmplitudes [2797] = 8'd114;
   assign soundFileAmplitudes [2798] = 8'd122;
   assign soundFileAmplitudes [2799] = 8'd131;
   assign soundFileAmplitudes [2800] = 8'd134;
   assign soundFileAmplitudes [2801] = 8'd127;
   assign soundFileAmplitudes [2802] = 8'd130;
   assign soundFileAmplitudes [2803] = 8'd138;
   assign soundFileAmplitudes [2804] = 8'd133;
   assign soundFileAmplitudes [2805] = 8'd146;
   assign soundFileAmplitudes [2806] = 8'd152;
   assign soundFileAmplitudes [2807] = 8'd146;
   assign soundFileAmplitudes [2808] = 8'd134;
   assign soundFileAmplitudes [2809] = 8'd110;
   assign soundFileAmplitudes [2810] = 8'd113;
   assign soundFileAmplitudes [2811] = 8'd106;
   assign soundFileAmplitudes [2812] = 8'd102;
   assign soundFileAmplitudes [2813] = 8'd90;
   assign soundFileAmplitudes [2814] = 8'd100;
   assign soundFileAmplitudes [2815] = 8'd112;
   assign soundFileAmplitudes [2816] = 8'd111;
   assign soundFileAmplitudes [2817] = 8'd107;
   assign soundFileAmplitudes [2818] = 8'd111;
   assign soundFileAmplitudes [2819] = 8'd119;
   assign soundFileAmplitudes [2820] = 8'd133;
   assign soundFileAmplitudes [2821] = 8'd131;
   assign soundFileAmplitudes [2822] = 8'd119;
   assign soundFileAmplitudes [2823] = 8'd110;
   assign soundFileAmplitudes [2824] = 8'd109;
   assign soundFileAmplitudes [2825] = 8'd115;
   assign soundFileAmplitudes [2826] = 8'd109;
   assign soundFileAmplitudes [2827] = 8'd130;
   assign soundFileAmplitudes [2828] = 8'd139;
   assign soundFileAmplitudes [2829] = 8'd139;
   assign soundFileAmplitudes [2830] = 8'd134;
   assign soundFileAmplitudes [2831] = 8'd135;
   assign soundFileAmplitudes [2832] = 8'd139;
   assign soundFileAmplitudes [2833] = 8'd143;
   assign soundFileAmplitudes [2834] = 8'd156;
   assign soundFileAmplitudes [2835] = 8'd161;
   assign soundFileAmplitudes [2836] = 8'd158;
   assign soundFileAmplitudes [2837] = 8'd159;
   assign soundFileAmplitudes [2838] = 8'd144;
   assign soundFileAmplitudes [2839] = 8'd144;
   assign soundFileAmplitudes [2840] = 8'd138;
   assign soundFileAmplitudes [2841] = 8'd114;
   assign soundFileAmplitudes [2842] = 8'd112;
   assign soundFileAmplitudes [2843] = 8'd115;
   assign soundFileAmplitudes [2844] = 8'd128;
   assign soundFileAmplitudes [2845] = 8'd128;
   assign soundFileAmplitudes [2846] = 8'd124;
   assign soundFileAmplitudes [2847] = 8'd113;
   assign soundFileAmplitudes [2848] = 8'd102;
   assign soundFileAmplitudes [2849] = 8'd100;
   assign soundFileAmplitudes [2850] = 8'd103;
   assign soundFileAmplitudes [2851] = 8'd105;
   assign soundFileAmplitudes [2852] = 8'd103;
   assign soundFileAmplitudes [2853] = 8'd110;
   assign soundFileAmplitudes [2854] = 8'd109;
   assign soundFileAmplitudes [2855] = 8'd95;
   assign soundFileAmplitudes [2856] = 8'd93;
   assign soundFileAmplitudes [2857] = 8'd110;
   assign soundFileAmplitudes [2858] = 8'd114;
   assign soundFileAmplitudes [2859] = 8'd114;
   assign soundFileAmplitudes [2860] = 8'd109;
   assign soundFileAmplitudes [2861] = 8'd116;
   assign soundFileAmplitudes [2862] = 8'd140;
   assign soundFileAmplitudes [2863] = 8'd146;
   assign soundFileAmplitudes [2864] = 8'd150;
   assign soundFileAmplitudes [2865] = 8'd156;
   assign soundFileAmplitudes [2866] = 8'd161;
   assign soundFileAmplitudes [2867] = 8'd159;
   assign soundFileAmplitudes [2868] = 8'd159;
   assign soundFileAmplitudes [2869] = 8'd154;
   assign soundFileAmplitudes [2870] = 8'd162;
   assign soundFileAmplitudes [2871] = 8'd156;
   assign soundFileAmplitudes [2872] = 8'd144;
   assign soundFileAmplitudes [2873] = 8'd149;
   assign soundFileAmplitudes [2874] = 8'd145;
   assign soundFileAmplitudes [2875] = 8'd142;
   assign soundFileAmplitudes [2876] = 8'd126;
   assign soundFileAmplitudes [2877] = 8'd128;
   assign soundFileAmplitudes [2878] = 8'd137;
   assign soundFileAmplitudes [2879] = 8'd141;
   assign soundFileAmplitudes [2880] = 8'd130;
   assign soundFileAmplitudes [2881] = 8'd115;
   assign soundFileAmplitudes [2882] = 8'd104;
   assign soundFileAmplitudes [2883] = 8'd100;
   assign soundFileAmplitudes [2884] = 8'd92;
   assign soundFileAmplitudes [2885] = 8'd87;
   assign soundFileAmplitudes [2886] = 8'd97;
   assign soundFileAmplitudes [2887] = 8'd91;
   assign soundFileAmplitudes [2888] = 8'd81;
   assign soundFileAmplitudes [2889] = 8'd88;
   assign soundFileAmplitudes [2890] = 8'd110;
   assign soundFileAmplitudes [2891] = 8'd130;
   assign soundFileAmplitudes [2892] = 8'd126;
   assign soundFileAmplitudes [2893] = 8'd117;
   assign soundFileAmplitudes [2894] = 8'd119;
   assign soundFileAmplitudes [2895] = 8'd129;
   assign soundFileAmplitudes [2896] = 8'd116;
   assign soundFileAmplitudes [2897] = 8'd104;
   assign soundFileAmplitudes [2898] = 8'd111;
   assign soundFileAmplitudes [2899] = 8'd123;
   assign soundFileAmplitudes [2900] = 8'd132;
   assign soundFileAmplitudes [2901] = 8'd136;
   assign soundFileAmplitudes [2902] = 8'd150;
   assign soundFileAmplitudes [2903] = 8'd133;
   assign soundFileAmplitudes [2904] = 8'd136;
   assign soundFileAmplitudes [2905] = 8'd133;
   assign soundFileAmplitudes [2906] = 8'd129;
   assign soundFileAmplitudes [2907] = 8'd154;
   assign soundFileAmplitudes [2908] = 8'd145;
   assign soundFileAmplitudes [2909] = 8'd145;
   assign soundFileAmplitudes [2910] = 8'd158;
   assign soundFileAmplitudes [2911] = 8'd161;
   assign soundFileAmplitudes [2912] = 8'd155;
   assign soundFileAmplitudes [2913] = 8'd135;
   assign soundFileAmplitudes [2914] = 8'd120;
   assign soundFileAmplitudes [2915] = 8'd127;
   assign soundFileAmplitudes [2916] = 8'd139;
   assign soundFileAmplitudes [2917] = 8'd131;
   assign soundFileAmplitudes [2918] = 8'd119;
   assign soundFileAmplitudes [2919] = 8'd109;
   assign soundFileAmplitudes [2920] = 8'd122;
   assign soundFileAmplitudes [2921] = 8'd137;
   assign soundFileAmplitudes [2922] = 8'd136;
   assign soundFileAmplitudes [2923] = 8'd133;
   assign soundFileAmplitudes [2924] = 8'd125;
   assign soundFileAmplitudes [2925] = 8'd113;
   assign soundFileAmplitudes [2926] = 8'd99;
   assign soundFileAmplitudes [2927] = 8'd110;
   assign soundFileAmplitudes [2928] = 8'd103;
   assign soundFileAmplitudes [2929] = 8'd90;
   assign soundFileAmplitudes [2930] = 8'd95;
   assign soundFileAmplitudes [2931] = 8'd113;
   assign soundFileAmplitudes [2932] = 8'd126;
   assign soundFileAmplitudes [2933] = 8'd118;
   assign soundFileAmplitudes [2934] = 8'd119;
   assign soundFileAmplitudes [2935] = 8'd117;
   assign soundFileAmplitudes [2936] = 8'd125;
   assign soundFileAmplitudes [2937] = 8'd128;
   assign soundFileAmplitudes [2938] = 8'd120;
   assign soundFileAmplitudes [2939] = 8'd128;
   assign soundFileAmplitudes [2940] = 8'd127;
   assign soundFileAmplitudes [2941] = 8'd137;
   assign soundFileAmplitudes [2942] = 8'd139;
   assign soundFileAmplitudes [2943] = 8'd129;
   assign soundFileAmplitudes [2944] = 8'd127;
   assign soundFileAmplitudes [2945] = 8'd133;
   assign soundFileAmplitudes [2946] = 8'd141;
   assign soundFileAmplitudes [2947] = 8'd141;
   assign soundFileAmplitudes [2948] = 8'd143;
   assign soundFileAmplitudes [2949] = 8'd152;
   assign soundFileAmplitudes [2950] = 8'd171;
   assign soundFileAmplitudes [2951] = 8'd159;
   assign soundFileAmplitudes [2952] = 8'd149;
   assign soundFileAmplitudes [2953] = 8'd154;
   assign soundFileAmplitudes [2954] = 8'd139;
   assign soundFileAmplitudes [2955] = 8'd122;
   assign soundFileAmplitudes [2956] = 8'd99;
   assign soundFileAmplitudes [2957] = 8'd95;
   assign soundFileAmplitudes [2958] = 8'd105;
   assign soundFileAmplitudes [2959] = 8'd89;
   assign soundFileAmplitudes [2960] = 8'd82;
   assign soundFileAmplitudes [2961] = 8'd94;
   assign soundFileAmplitudes [2962] = 8'd108;
   assign soundFileAmplitudes [2963] = 8'd112;
   assign soundFileAmplitudes [2964] = 8'd121;
   assign soundFileAmplitudes [2965] = 8'd115;
   assign soundFileAmplitudes [2966] = 8'd129;
   assign soundFileAmplitudes [2967] = 8'd128;
   assign soundFileAmplitudes [2968] = 8'd121;
   assign soundFileAmplitudes [2969] = 8'd113;
   assign soundFileAmplitudes [2970] = 8'd104;
   assign soundFileAmplitudes [2971] = 8'd113;
   assign soundFileAmplitudes [2972] = 8'd99;
   assign soundFileAmplitudes [2973] = 8'd117;
   assign soundFileAmplitudes [2974] = 8'd121;
   assign soundFileAmplitudes [2975] = 8'd124;
   assign soundFileAmplitudes [2976] = 8'd118;
   assign soundFileAmplitudes [2977] = 8'd115;
   assign soundFileAmplitudes [2978] = 8'd146;
   assign soundFileAmplitudes [2979] = 8'd163;
   assign soundFileAmplitudes [2980] = 8'd176;
   assign soundFileAmplitudes [2981] = 8'd177;
   assign soundFileAmplitudes [2982] = 8'd164;
   assign soundFileAmplitudes [2983] = 8'd172;
   assign soundFileAmplitudes [2984] = 8'd153;
   assign soundFileAmplitudes [2985] = 8'd143;
   assign soundFileAmplitudes [2986] = 8'd156;
   assign soundFileAmplitudes [2987] = 8'd126;
   assign soundFileAmplitudes [2988] = 8'd104;
   assign soundFileAmplitudes [2989] = 8'd104;
   assign soundFileAmplitudes [2990] = 8'd116;
   assign soundFileAmplitudes [2991] = 8'd113;
   assign soundFileAmplitudes [2992] = 8'd101;
   assign soundFileAmplitudes [2993] = 8'd95;
   assign soundFileAmplitudes [2994] = 8'd99;
   assign soundFileAmplitudes [2995] = 8'd124;
   assign soundFileAmplitudes [2996] = 8'd128;
   assign soundFileAmplitudes [2997] = 8'd142;
   assign soundFileAmplitudes [2998] = 8'd135;
   assign soundFileAmplitudes [2999] = 8'd128;
   assign soundFileAmplitudes [3000] = 8'd122;
   assign soundFileAmplitudes [3001] = 8'd94;
   assign soundFileAmplitudes [3002] = 8'd106;
   assign soundFileAmplitudes [3003] = 8'd110;
   assign soundFileAmplitudes [3004] = 8'd121;
   assign soundFileAmplitudes [3005] = 8'd109;
   assign soundFileAmplitudes [3006] = 8'd101;
   assign soundFileAmplitudes [3007] = 8'd105;
   assign soundFileAmplitudes [3008] = 8'd120;
   assign soundFileAmplitudes [3009] = 8'd139;
   assign soundFileAmplitudes [3010] = 8'd130;
   assign soundFileAmplitudes [3011] = 8'd137;
   assign soundFileAmplitudes [3012] = 8'd150;
   assign soundFileAmplitudes [3013] = 8'd137;
   assign soundFileAmplitudes [3014] = 8'd140;
   assign soundFileAmplitudes [3015] = 8'd158;
   assign soundFileAmplitudes [3016] = 8'd143;
   assign soundFileAmplitudes [3017] = 8'd144;
   assign soundFileAmplitudes [3018] = 8'd131;
   assign soundFileAmplitudes [3019] = 8'd130;
   assign soundFileAmplitudes [3020] = 8'd144;
   assign soundFileAmplitudes [3021] = 8'd141;
   assign soundFileAmplitudes [3022] = 8'd146;
   assign soundFileAmplitudes [3023] = 8'd137;
   assign soundFileAmplitudes [3024] = 8'd122;
   assign soundFileAmplitudes [3025] = 8'd130;
   assign soundFileAmplitudes [3026] = 8'd137;
   assign soundFileAmplitudes [3027] = 8'd129;
   assign soundFileAmplitudes [3028] = 8'd99;
   assign soundFileAmplitudes [3029] = 8'd78;
   assign soundFileAmplitudes [3030] = 8'd68;
   assign soundFileAmplitudes [3031] = 8'd86;
   assign soundFileAmplitudes [3032] = 8'd112;
   assign soundFileAmplitudes [3033] = 8'd117;
   assign soundFileAmplitudes [3034] = 8'd134;
   assign soundFileAmplitudes [3035] = 8'd137;
   assign soundFileAmplitudes [3036] = 8'd142;
   assign soundFileAmplitudes [3037] = 8'd155;
   assign soundFileAmplitudes [3038] = 8'd154;
   assign soundFileAmplitudes [3039] = 8'd138;
   assign soundFileAmplitudes [3040] = 8'd122;
   assign soundFileAmplitudes [3041] = 8'd117;
   assign soundFileAmplitudes [3042] = 8'd119;
   assign soundFileAmplitudes [3043] = 8'd122;
   assign soundFileAmplitudes [3044] = 8'd123;
   assign soundFileAmplitudes [3045] = 8'd107;
   assign soundFileAmplitudes [3046] = 8'd106;
   assign soundFileAmplitudes [3047] = 8'd111;
   assign soundFileAmplitudes [3048] = 8'd117;
   assign soundFileAmplitudes [3049] = 8'd128;
   assign soundFileAmplitudes [3050] = 8'd133;
   assign soundFileAmplitudes [3051] = 8'd140;
   assign soundFileAmplitudes [3052] = 8'd151;
   assign soundFileAmplitudes [3053] = 8'd151;
   assign soundFileAmplitudes [3054] = 8'd148;
   assign soundFileAmplitudes [3055] = 8'd142;
   assign soundFileAmplitudes [3056] = 8'd135;
   assign soundFileAmplitudes [3057] = 8'd149;
   assign soundFileAmplitudes [3058] = 8'd147;
   assign soundFileAmplitudes [3059] = 8'd143;
   assign soundFileAmplitudes [3060] = 8'd113;
   assign soundFileAmplitudes [3061] = 8'd94;
   assign soundFileAmplitudes [3062] = 8'd88;
   assign soundFileAmplitudes [3063] = 8'd112;
   assign soundFileAmplitudes [3064] = 8'd116;
   assign soundFileAmplitudes [3065] = 8'd100;
   assign soundFileAmplitudes [3066] = 8'd115;
   assign soundFileAmplitudes [3067] = 8'd106;
   assign soundFileAmplitudes [3068] = 8'd122;
   assign soundFileAmplitudes [3069] = 8'd132;
   assign soundFileAmplitudes [3070] = 8'd136;
   assign soundFileAmplitudes [3071] = 8'd145;
   assign soundFileAmplitudes [3072] = 8'd137;
   assign soundFileAmplitudes [3073] = 8'd124;
   assign soundFileAmplitudes [3074] = 8'd129;
   assign soundFileAmplitudes [3075] = 8'd137;
   assign soundFileAmplitudes [3076] = 8'd121;
   assign soundFileAmplitudes [3077] = 8'd105;
   assign soundFileAmplitudes [3078] = 8'd119;
   assign soundFileAmplitudes [3079] = 8'd125;
   assign soundFileAmplitudes [3080] = 8'd125;
   assign soundFileAmplitudes [3081] = 8'd117;
   assign soundFileAmplitudes [3082] = 8'd110;
   assign soundFileAmplitudes [3083] = 8'd119;
   assign soundFileAmplitudes [3084] = 8'd133;
   assign soundFileAmplitudes [3085] = 8'd125;
   assign soundFileAmplitudes [3086] = 8'd133;
   assign soundFileAmplitudes [3087] = 8'd140;
   assign soundFileAmplitudes [3088] = 8'd111;
   assign soundFileAmplitudes [3089] = 8'd120;
   assign soundFileAmplitudes [3090] = 8'd123;
   assign soundFileAmplitudes [3091] = 8'd136;
   assign soundFileAmplitudes [3092] = 8'd139;
   assign soundFileAmplitudes [3093] = 8'd140;
   assign soundFileAmplitudes [3094] = 8'd147;
   assign soundFileAmplitudes [3095] = 8'd148;
   assign soundFileAmplitudes [3096] = 8'd151;
   assign soundFileAmplitudes [3097] = 8'd143;
   assign soundFileAmplitudes [3098] = 8'd138;
   assign soundFileAmplitudes [3099] = 8'd129;
   assign soundFileAmplitudes [3100] = 8'd135;
   assign soundFileAmplitudes [3101] = 8'd122;
   assign soundFileAmplitudes [3102] = 8'd109;
   assign soundFileAmplitudes [3103] = 8'd101;
   assign soundFileAmplitudes [3104] = 8'd92;
   assign soundFileAmplitudes [3105] = 8'd97;
   assign soundFileAmplitudes [3106] = 8'd108;
   assign soundFileAmplitudes [3107] = 8'd128;
   assign soundFileAmplitudes [3108] = 8'd127;
   assign soundFileAmplitudes [3109] = 8'd132;
   assign soundFileAmplitudes [3110] = 8'd125;
   assign soundFileAmplitudes [3111] = 8'd113;
   assign soundFileAmplitudes [3112] = 8'd113;
   assign soundFileAmplitudes [3113] = 8'd111;
   assign soundFileAmplitudes [3114] = 8'd132;
   assign soundFileAmplitudes [3115] = 8'd134;
   assign soundFileAmplitudes [3116] = 8'd125;
   assign soundFileAmplitudes [3117] = 8'd125;
   assign soundFileAmplitudes [3118] = 8'd119;
   assign soundFileAmplitudes [3119] = 8'd103;
   assign soundFileAmplitudes [3120] = 8'd106;
   assign soundFileAmplitudes [3121] = 8'd116;
   assign soundFileAmplitudes [3122] = 8'd128;
   assign soundFileAmplitudes [3123] = 8'd134;
   assign soundFileAmplitudes [3124] = 8'd128;
   assign soundFileAmplitudes [3125] = 8'd133;
   assign soundFileAmplitudes [3126] = 8'd141;
   assign soundFileAmplitudes [3127] = 8'd147;
   assign soundFileAmplitudes [3128] = 8'd156;
   assign soundFileAmplitudes [3129] = 8'd162;
   assign soundFileAmplitudes [3130] = 8'd163;
   assign soundFileAmplitudes [3131] = 8'd162;
   assign soundFileAmplitudes [3132] = 8'd155;
   assign soundFileAmplitudes [3133] = 8'd140;
   assign soundFileAmplitudes [3134] = 8'd115;
   assign soundFileAmplitudes [3135] = 8'd101;
   assign soundFileAmplitudes [3136] = 8'd100;
   assign soundFileAmplitudes [3137] = 8'd110;
   assign soundFileAmplitudes [3138] = 8'd111;
   assign soundFileAmplitudes [3139] = 8'd99;
   assign soundFileAmplitudes [3140] = 8'd95;
   assign soundFileAmplitudes [3141] = 8'd87;
   assign soundFileAmplitudes [3142] = 8'd97;
   assign soundFileAmplitudes [3143] = 8'd113;
   assign soundFileAmplitudes [3144] = 8'd120;
   assign soundFileAmplitudes [3145] = 8'd134;
   assign soundFileAmplitudes [3146] = 8'd147;
   assign soundFileAmplitudes [3147] = 8'd143;
   assign soundFileAmplitudes [3148] = 8'd139;
   assign soundFileAmplitudes [3149] = 8'd140;
   assign soundFileAmplitudes [3150] = 8'd126;
   assign soundFileAmplitudes [3151] = 8'd128;
   assign soundFileAmplitudes [3152] = 8'd121;
   assign soundFileAmplitudes [3153] = 8'd114;
   assign soundFileAmplitudes [3154] = 8'd116;
   assign soundFileAmplitudes [3155] = 8'd105;
   assign soundFileAmplitudes [3156] = 8'd118;
   assign soundFileAmplitudes [3157] = 8'd122;
   assign soundFileAmplitudes [3158] = 8'd132;
   assign soundFileAmplitudes [3159] = 8'd148;
   assign soundFileAmplitudes [3160] = 8'd149;
   assign soundFileAmplitudes [3161] = 8'd139;
   assign soundFileAmplitudes [3162] = 8'd135;
   assign soundFileAmplitudes [3163] = 8'd140;
   assign soundFileAmplitudes [3164] = 8'd140;
   assign soundFileAmplitudes [3165] = 8'd151;
   assign soundFileAmplitudes [3166] = 8'd142;
   assign soundFileAmplitudes [3167] = 8'd140;
   assign soundFileAmplitudes [3168] = 8'd142;
   assign soundFileAmplitudes [3169] = 8'd136;
   assign soundFileAmplitudes [3170] = 8'd121;
   assign soundFileAmplitudes [3171] = 8'd113;
   assign soundFileAmplitudes [3172] = 8'd111;
   assign soundFileAmplitudes [3173] = 8'd102;
   assign soundFileAmplitudes [3174] = 8'd110;
   assign soundFileAmplitudes [3175] = 8'd104;
   assign soundFileAmplitudes [3176] = 8'd101;
   assign soundFileAmplitudes [3177] = 8'd110;
   assign soundFileAmplitudes [3178] = 8'd113;
   assign soundFileAmplitudes [3179] = 8'd128;
   assign soundFileAmplitudes [3180] = 8'd118;
   assign soundFileAmplitudes [3181] = 8'd114;
   assign soundFileAmplitudes [3182] = 8'd118;
   assign soundFileAmplitudes [3183] = 8'd117;
   assign soundFileAmplitudes [3184] = 8'd135;
   assign soundFileAmplitudes [3185] = 8'd140;
   assign soundFileAmplitudes [3186] = 8'd135;
   assign soundFileAmplitudes [3187] = 8'd143;
   assign soundFileAmplitudes [3188] = 8'd146;
   assign soundFileAmplitudes [3189] = 8'd135;
   assign soundFileAmplitudes [3190] = 8'd126;
   assign soundFileAmplitudes [3191] = 8'd130;
   assign soundFileAmplitudes [3192] = 8'd138;
   assign soundFileAmplitudes [3193] = 8'd128;
   assign soundFileAmplitudes [3194] = 8'd120;
   assign soundFileAmplitudes [3195] = 8'd113;
   assign soundFileAmplitudes [3196] = 8'd117;
   assign soundFileAmplitudes [3197] = 8'd114;
   assign soundFileAmplitudes [3198] = 8'd118;
   assign soundFileAmplitudes [3199] = 8'd122;
   assign soundFileAmplitudes [3200] = 8'd129;
   assign soundFileAmplitudes [3201] = 8'd132;
   assign soundFileAmplitudes [3202] = 8'd136;
   assign soundFileAmplitudes [3203] = 8'd155;
   assign soundFileAmplitudes [3204] = 8'd141;
   assign soundFileAmplitudes [3205] = 8'd135;
   assign soundFileAmplitudes [3206] = 8'd123;
   assign soundFileAmplitudes [3207] = 8'd119;
   assign soundFileAmplitudes [3208] = 8'd130;
   assign soundFileAmplitudes [3209] = 8'd131;
   assign soundFileAmplitudes [3210] = 8'd132;
   assign soundFileAmplitudes [3211] = 8'd107;
   assign soundFileAmplitudes [3212] = 8'd96;
   assign soundFileAmplitudes [3213] = 8'd112;
   assign soundFileAmplitudes [3214] = 8'd105;
   assign soundFileAmplitudes [3215] = 8'd104;
   assign soundFileAmplitudes [3216] = 8'd112;
   assign soundFileAmplitudes [3217] = 8'd126;
   assign soundFileAmplitudes [3218] = 8'd128;
   assign soundFileAmplitudes [3219] = 8'd126;
   assign soundFileAmplitudes [3220] = 8'd133;
   assign soundFileAmplitudes [3221] = 8'd130;
   assign soundFileAmplitudes [3222] = 8'd123;
   assign soundFileAmplitudes [3223] = 8'd133;
   assign soundFileAmplitudes [3224] = 8'd146;
   assign soundFileAmplitudes [3225] = 8'd134;
   assign soundFileAmplitudes [3226] = 8'd136;
   assign soundFileAmplitudes [3227] = 8'd131;
   assign soundFileAmplitudes [3228] = 8'd137;
   assign soundFileAmplitudes [3229] = 8'd137;
   assign soundFileAmplitudes [3230] = 8'd133;
   assign soundFileAmplitudes [3231] = 8'd128;
   assign soundFileAmplitudes [3232] = 8'd124;
   assign soundFileAmplitudes [3233] = 8'd120;
   assign soundFileAmplitudes [3234] = 8'd119;
   assign soundFileAmplitudes [3235] = 8'd131;
   assign soundFileAmplitudes [3236] = 8'd134;
   assign soundFileAmplitudes [3237] = 8'd131;
   assign soundFileAmplitudes [3238] = 8'd114;
   assign soundFileAmplitudes [3239] = 8'd111;
   assign soundFileAmplitudes [3240] = 8'd94;
   assign soundFileAmplitudes [3241] = 8'd107;
   assign soundFileAmplitudes [3242] = 8'd125;
   assign soundFileAmplitudes [3243] = 8'd115;
   assign soundFileAmplitudes [3244] = 8'd106;
   assign soundFileAmplitudes [3245] = 8'd103;
   assign soundFileAmplitudes [3246] = 8'd115;
   assign soundFileAmplitudes [3247] = 8'd127;
   assign soundFileAmplitudes [3248] = 8'd136;
   assign soundFileAmplitudes [3249] = 8'd138;
   assign soundFileAmplitudes [3250] = 8'd135;
   assign soundFileAmplitudes [3251] = 8'd135;
   assign soundFileAmplitudes [3252] = 8'd129;
   assign soundFileAmplitudes [3253] = 8'd116;
   assign soundFileAmplitudes [3254] = 8'd129;
   assign soundFileAmplitudes [3255] = 8'd137;
   assign soundFileAmplitudes [3256] = 8'd124;
   assign soundFileAmplitudes [3257] = 8'd123;
   assign soundFileAmplitudes [3258] = 8'd128;
   assign soundFileAmplitudes [3259] = 8'd139;
   assign soundFileAmplitudes [3260] = 8'd140;
   assign soundFileAmplitudes [3261] = 8'd135;
   assign soundFileAmplitudes [3262] = 8'd149;
   assign soundFileAmplitudes [3263] = 8'd156;
   assign soundFileAmplitudes [3264] = 8'd151;
   assign soundFileAmplitudes [3265] = 8'd157;
   assign soundFileAmplitudes [3266] = 8'd145;
   assign soundFileAmplitudes [3267] = 8'd129;
   assign soundFileAmplitudes [3268] = 8'd118;
   assign soundFileAmplitudes [3269] = 8'd97;
   assign soundFileAmplitudes [3270] = 8'd96;
   assign soundFileAmplitudes [3271] = 8'd100;
   assign soundFileAmplitudes [3272] = 8'd104;
   assign soundFileAmplitudes [3273] = 8'd107;
   assign soundFileAmplitudes [3274] = 8'd105;
   assign soundFileAmplitudes [3275] = 8'd109;
   assign soundFileAmplitudes [3276] = 8'd116;
   assign soundFileAmplitudes [3277] = 8'd128;
   assign soundFileAmplitudes [3278] = 8'd127;
   assign soundFileAmplitudes [3279] = 8'd136;
   assign soundFileAmplitudes [3280] = 8'd153;
   assign soundFileAmplitudes [3281] = 8'd145;
   assign soundFileAmplitudes [3282] = 8'd129;
   assign soundFileAmplitudes [3283] = 8'd124;
   assign soundFileAmplitudes [3284] = 8'd123;
   assign soundFileAmplitudes [3285] = 8'd123;
   assign soundFileAmplitudes [3286] = 8'd105;
   assign soundFileAmplitudes [3287] = 8'd106;
   assign soundFileAmplitudes [3288] = 8'd118;
   assign soundFileAmplitudes [3289] = 8'd115;
   assign soundFileAmplitudes [3290] = 8'd124;
   assign soundFileAmplitudes [3291] = 8'd125;
   assign soundFileAmplitudes [3292] = 8'd129;
   assign soundFileAmplitudes [3293] = 8'd122;
   assign soundFileAmplitudes [3294] = 8'd129;
   assign soundFileAmplitudes [3295] = 8'd152;
   assign soundFileAmplitudes [3296] = 8'd143;
   assign soundFileAmplitudes [3297] = 8'd136;
   assign soundFileAmplitudes [3298] = 8'd132;
   assign soundFileAmplitudes [3299] = 8'd113;
   assign soundFileAmplitudes [3300] = 8'd114;
   assign soundFileAmplitudes [3301] = 8'd127;
   assign soundFileAmplitudes [3302] = 8'd115;
   assign soundFileAmplitudes [3303] = 8'd121;
   assign soundFileAmplitudes [3304] = 8'd123;
   assign soundFileAmplitudes [3305] = 8'd133;
   assign soundFileAmplitudes [3306] = 8'd156;
   assign soundFileAmplitudes [3307] = 8'd160;
   assign soundFileAmplitudes [3308] = 8'd145;
   assign soundFileAmplitudes [3309] = 8'd146;
   assign soundFileAmplitudes [3310] = 8'd149;
   assign soundFileAmplitudes [3311] = 8'd131;
   assign soundFileAmplitudes [3312] = 8'd124;
   assign soundFileAmplitudes [3313] = 8'd120;
   assign soundFileAmplitudes [3314] = 8'd118;
   assign soundFileAmplitudes [3315] = 8'd110;
   assign soundFileAmplitudes [3316] = 8'd114;
   assign soundFileAmplitudes [3317] = 8'd120;
   assign soundFileAmplitudes [3318] = 8'd128;
   assign soundFileAmplitudes [3319] = 8'd121;
   assign soundFileAmplitudes [3320] = 8'd116;
   assign soundFileAmplitudes [3321] = 8'd119;
   assign soundFileAmplitudes [3322] = 8'd137;
   assign soundFileAmplitudes [3323] = 8'd133;
   assign soundFileAmplitudes [3324] = 8'd124;
   assign soundFileAmplitudes [3325] = 8'd113;
   assign soundFileAmplitudes [3326] = 8'd94;
   assign soundFileAmplitudes [3327] = 8'd97;
   assign soundFileAmplitudes [3328] = 8'd82;
   assign soundFileAmplitudes [3329] = 8'd91;
   assign soundFileAmplitudes [3330] = 8'd99;
   assign soundFileAmplitudes [3331] = 8'd100;
   assign soundFileAmplitudes [3332] = 8'd118;
   assign soundFileAmplitudes [3333] = 8'd129;
   assign soundFileAmplitudes [3334] = 8'd141;
   assign soundFileAmplitudes [3335] = 8'd160;
   assign soundFileAmplitudes [3336] = 8'd165;
   assign soundFileAmplitudes [3337] = 8'd161;
   assign soundFileAmplitudes [3338] = 8'd157;
   assign soundFileAmplitudes [3339] = 8'd159;
   assign soundFileAmplitudes [3340] = 8'd158;
   assign soundFileAmplitudes [3341] = 8'd158;
   assign soundFileAmplitudes [3342] = 8'd150;
   assign soundFileAmplitudes [3343] = 8'd137;
   assign soundFileAmplitudes [3344] = 8'd113;
   assign soundFileAmplitudes [3345] = 8'd103;
   assign soundFileAmplitudes [3346] = 8'd100;
   assign soundFileAmplitudes [3347] = 8'd110;
   assign soundFileAmplitudes [3348] = 8'd120;
   assign soundFileAmplitudes [3349] = 8'd113;
   assign soundFileAmplitudes [3350] = 8'd113;
   assign soundFileAmplitudes [3351] = 8'd117;
   assign soundFileAmplitudes [3352] = 8'd122;
   assign soundFileAmplitudes [3353] = 8'd132;
   assign soundFileAmplitudes [3354] = 8'd144;
   assign soundFileAmplitudes [3355] = 8'd115;
   assign soundFileAmplitudes [3356] = 8'd114;
   assign soundFileAmplitudes [3357] = 8'd101;
   assign soundFileAmplitudes [3358] = 8'd101;
   assign soundFileAmplitudes [3359] = 8'd103;
   assign soundFileAmplitudes [3360] = 8'd88;
   assign soundFileAmplitudes [3361] = 8'd97;
   assign soundFileAmplitudes [3362] = 8'd101;
   assign soundFileAmplitudes [3363] = 8'd108;
   assign soundFileAmplitudes [3364] = 8'd129;
   assign soundFileAmplitudes [3365] = 8'd135;
   assign soundFileAmplitudes [3366] = 8'd137;
   assign soundFileAmplitudes [3367] = 8'd141;
   assign soundFileAmplitudes [3368] = 8'd147;
   assign soundFileAmplitudes [3369] = 8'd163;
   assign soundFileAmplitudes [3370] = 8'd164;
   assign soundFileAmplitudes [3371] = 8'd163;
   assign soundFileAmplitudes [3372] = 8'd163;
   assign soundFileAmplitudes [3373] = 8'd152;
   assign soundFileAmplitudes [3374] = 8'd133;
   assign soundFileAmplitudes [3375] = 8'd118;
   assign soundFileAmplitudes [3376] = 8'd127;
   assign soundFileAmplitudes [3377] = 8'd148;
   assign soundFileAmplitudes [3378] = 8'd139;
   assign soundFileAmplitudes [3379] = 8'd141;
   assign soundFileAmplitudes [3380] = 8'd131;
   assign soundFileAmplitudes [3381] = 8'd130;
   assign soundFileAmplitudes [3382] = 8'd112;
   assign soundFileAmplitudes [3383] = 8'd121;
   assign soundFileAmplitudes [3384] = 8'd126;
   assign soundFileAmplitudes [3385] = 8'd106;
   assign soundFileAmplitudes [3386] = 8'd104;
   assign soundFileAmplitudes [3387] = 8'd82;
   assign soundFileAmplitudes [3388] = 8'd100;
   assign soundFileAmplitudes [3389] = 8'd107;
   assign soundFileAmplitudes [3390] = 8'd116;
   assign soundFileAmplitudes [3391] = 8'd110;
   assign soundFileAmplitudes [3392] = 8'd96;
   assign soundFileAmplitudes [3393] = 8'd104;
   assign soundFileAmplitudes [3394] = 8'd120;
   assign soundFileAmplitudes [3395] = 8'd136;
   assign soundFileAmplitudes [3396] = 8'd137;
   assign soundFileAmplitudes [3397] = 8'd123;
   assign soundFileAmplitudes [3398] = 8'd125;
   assign soundFileAmplitudes [3399] = 8'd142;
   assign soundFileAmplitudes [3400] = 8'd146;
   assign soundFileAmplitudes [3401] = 8'd144;
   assign soundFileAmplitudes [3402] = 8'd136;
   assign soundFileAmplitudes [3403] = 8'd114;
   assign soundFileAmplitudes [3404] = 8'd108;
   assign soundFileAmplitudes [3405] = 8'd129;
   assign soundFileAmplitudes [3406] = 8'd140;
   assign soundFileAmplitudes [3407] = 8'd145;
   assign soundFileAmplitudes [3408] = 8'd129;
   assign soundFileAmplitudes [3409] = 8'd125;
   assign soundFileAmplitudes [3410] = 8'd133;
   assign soundFileAmplitudes [3411] = 8'd135;
   assign soundFileAmplitudes [3412] = 8'd126;
   assign soundFileAmplitudes [3413] = 8'd143;
   assign soundFileAmplitudes [3414] = 8'd151;
   assign soundFileAmplitudes [3415] = 8'd137;
   assign soundFileAmplitudes [3416] = 8'd121;
   assign soundFileAmplitudes [3417] = 8'd95;
   assign soundFileAmplitudes [3418] = 8'd105;
   assign soundFileAmplitudes [3419] = 8'd98;
   assign soundFileAmplitudes [3420] = 8'd103;
   assign soundFileAmplitudes [3421] = 8'd111;
   assign soundFileAmplitudes [3422] = 8'd107;
   assign soundFileAmplitudes [3423] = 8'd111;
   assign soundFileAmplitudes [3424] = 8'd114;
   assign soundFileAmplitudes [3425] = 8'd131;
   assign soundFileAmplitudes [3426] = 8'd147;
   assign soundFileAmplitudes [3427] = 8'd155;
   assign soundFileAmplitudes [3428] = 8'd156;
   assign soundFileAmplitudes [3429] = 8'd141;
   assign soundFileAmplitudes [3430] = 8'd129;
   assign soundFileAmplitudes [3431] = 8'd141;
   assign soundFileAmplitudes [3432] = 8'd137;
   assign soundFileAmplitudes [3433] = 8'd124;
   assign soundFileAmplitudes [3434] = 8'd109;
   assign soundFileAmplitudes [3435] = 8'd115;
   assign soundFileAmplitudes [3436] = 8'd133;
   assign soundFileAmplitudes [3437] = 8'd146;
   assign soundFileAmplitudes [3438] = 8'd134;
   assign soundFileAmplitudes [3439] = 8'd117;
   assign soundFileAmplitudes [3440] = 8'd106;
   assign soundFileAmplitudes [3441] = 8'd126;
   assign soundFileAmplitudes [3442] = 8'd123;
   assign soundFileAmplitudes [3443] = 8'd122;
   assign soundFileAmplitudes [3444] = 8'd138;
   assign soundFileAmplitudes [3445] = 8'd111;
   assign soundFileAmplitudes [3446] = 8'd115;
   assign soundFileAmplitudes [3447] = 8'd83;
   assign soundFileAmplitudes [3448] = 8'd83;
   assign soundFileAmplitudes [3449] = 8'd114;
   assign soundFileAmplitudes [3450] = 8'd123;
   assign soundFileAmplitudes [3451] = 8'd124;
   assign soundFileAmplitudes [3452] = 8'd120;
   assign soundFileAmplitudes [3453] = 8'd130;
   assign soundFileAmplitudes [3454] = 8'd142;
   assign soundFileAmplitudes [3455] = 8'd153;
   assign soundFileAmplitudes [3456] = 8'd160;
   assign soundFileAmplitudes [3457] = 8'd171;
   assign soundFileAmplitudes [3458] = 8'd158;
   assign soundFileAmplitudes [3459] = 8'd150;
   assign soundFileAmplitudes [3460] = 8'd142;
   assign soundFileAmplitudes [3461] = 8'd132;
   assign soundFileAmplitudes [3462] = 8'd130;
   assign soundFileAmplitudes [3463] = 8'd123;
   assign soundFileAmplitudes [3464] = 8'd117;
   assign soundFileAmplitudes [3465] = 8'd119;
   assign soundFileAmplitudes [3466] = 8'd125;
   assign soundFileAmplitudes [3467] = 8'd127;
   assign soundFileAmplitudes [3468] = 8'd120;
   assign soundFileAmplitudes [3469] = 8'd111;
   assign soundFileAmplitudes [3470] = 8'd108;
   assign soundFileAmplitudes [3471] = 8'd123;
   assign soundFileAmplitudes [3472] = 8'd129;
   assign soundFileAmplitudes [3473] = 8'd124;
   assign soundFileAmplitudes [3474] = 8'd123;
   assign soundFileAmplitudes [3475] = 8'd110;
   assign soundFileAmplitudes [3476] = 8'd108;
   assign soundFileAmplitudes [3477] = 8'd97;
   assign soundFileAmplitudes [3478] = 8'd81;
   assign soundFileAmplitudes [3479] = 8'd104;
   assign soundFileAmplitudes [3480] = 8'd113;
   assign soundFileAmplitudes [3481] = 8'd104;
   assign soundFileAmplitudes [3482] = 8'd110;
   assign soundFileAmplitudes [3483] = 8'd104;
   assign soundFileAmplitudes [3484] = 8'd111;
   assign soundFileAmplitudes [3485] = 8'd133;
   assign soundFileAmplitudes [3486] = 8'd157;
   assign soundFileAmplitudes [3487] = 8'd172;
   assign soundFileAmplitudes [3488] = 8'd165;
   assign soundFileAmplitudes [3489] = 8'd157;
   assign soundFileAmplitudes [3490] = 8'd143;
   assign soundFileAmplitudes [3491] = 8'd141;
   assign soundFileAmplitudes [3492] = 8'd140;
   assign soundFileAmplitudes [3493] = 8'd133;
   assign soundFileAmplitudes [3494] = 8'd130;
   assign soundFileAmplitudes [3495] = 8'd127;
   assign soundFileAmplitudes [3496] = 8'd132;
   assign soundFileAmplitudes [3497] = 8'd138;
   assign soundFileAmplitudes [3498] = 8'd132;
   assign soundFileAmplitudes [3499] = 8'd113;
   assign soundFileAmplitudes [3500] = 8'd108;
   assign soundFileAmplitudes [3501] = 8'd120;
   assign soundFileAmplitudes [3502] = 8'd138;
   assign soundFileAmplitudes [3503] = 8'd134;
   assign soundFileAmplitudes [3504] = 8'd133;
   assign soundFileAmplitudes [3505] = 8'd121;
   assign soundFileAmplitudes [3506] = 8'd112;
   assign soundFileAmplitudes [3507] = 8'd95;
   assign soundFileAmplitudes [3508] = 8'd87;
   assign soundFileAmplitudes [3509] = 8'd107;
   assign soundFileAmplitudes [3510] = 8'd105;
   assign soundFileAmplitudes [3511] = 8'd104;
   assign soundFileAmplitudes [3512] = 8'd91;
   assign soundFileAmplitudes [3513] = 8'd102;
   assign soundFileAmplitudes [3514] = 8'd119;
   assign soundFileAmplitudes [3515] = 8'd137;
   assign soundFileAmplitudes [3516] = 8'd142;
   assign soundFileAmplitudes [3517] = 8'd134;
   assign soundFileAmplitudes [3518] = 8'd145;
   assign soundFileAmplitudes [3519] = 8'd148;
   assign soundFileAmplitudes [3520] = 8'd145;
   assign soundFileAmplitudes [3521] = 8'd139;
   assign soundFileAmplitudes [3522] = 8'd148;
   assign soundFileAmplitudes [3523] = 8'd144;
   assign soundFileAmplitudes [3524] = 8'd137;
   assign soundFileAmplitudes [3525] = 8'd126;
   assign soundFileAmplitudes [3526] = 8'd121;
   assign soundFileAmplitudes [3527] = 8'd137;
   assign soundFileAmplitudes [3528] = 8'd152;
   assign soundFileAmplitudes [3529] = 8'd143;
   assign soundFileAmplitudes [3530] = 8'd124;
   assign soundFileAmplitudes [3531] = 8'd121;
   assign soundFileAmplitudes [3532] = 8'd132;
   assign soundFileAmplitudes [3533] = 8'd141;
   assign soundFileAmplitudes [3534] = 8'd146;
   assign soundFileAmplitudes [3535] = 8'd137;
   assign soundFileAmplitudes [3536] = 8'd113;
   assign soundFileAmplitudes [3537] = 8'd109;
   assign soundFileAmplitudes [3538] = 8'd98;
   assign soundFileAmplitudes [3539] = 8'd99;
   assign soundFileAmplitudes [3540] = 8'd108;
   assign soundFileAmplitudes [3541] = 8'd99;
   assign soundFileAmplitudes [3542] = 8'd103;
   assign soundFileAmplitudes [3543] = 8'd108;
   assign soundFileAmplitudes [3544] = 8'd117;
   assign soundFileAmplitudes [3545] = 8'd126;
   assign soundFileAmplitudes [3546] = 8'd128;
   assign soundFileAmplitudes [3547] = 8'd133;
   assign soundFileAmplitudes [3548] = 8'd133;
   assign soundFileAmplitudes [3549] = 8'd152;
   assign soundFileAmplitudes [3550] = 8'd147;
   assign soundFileAmplitudes [3551] = 8'd135;
   assign soundFileAmplitudes [3552] = 8'd127;
   assign soundFileAmplitudes [3553] = 8'd112;
   assign soundFileAmplitudes [3554] = 8'd117;
   assign soundFileAmplitudes [3555] = 8'd106;
   assign soundFileAmplitudes [3556] = 8'd101;
   assign soundFileAmplitudes [3557] = 8'd121;
   assign soundFileAmplitudes [3558] = 8'd127;
   assign soundFileAmplitudes [3559] = 8'd122;
   assign soundFileAmplitudes [3560] = 8'd128;
   assign soundFileAmplitudes [3561] = 8'd129;
   assign soundFileAmplitudes [3562] = 8'd134;
   assign soundFileAmplitudes [3563] = 8'd132;
   assign soundFileAmplitudes [3564] = 8'd126;
   assign soundFileAmplitudes [3565] = 8'd139;
   assign soundFileAmplitudes [3566] = 8'd147;
   assign soundFileAmplitudes [3567] = 8'd144;
   assign soundFileAmplitudes [3568] = 8'd122;
   assign soundFileAmplitudes [3569] = 8'd107;
   assign soundFileAmplitudes [3570] = 8'd115;
   assign soundFileAmplitudes [3571] = 8'd125;
   assign soundFileAmplitudes [3572] = 8'd122;
   assign soundFileAmplitudes [3573] = 8'd111;
   assign soundFileAmplitudes [3574] = 8'd103;
   assign soundFileAmplitudes [3575] = 8'd130;
   assign soundFileAmplitudes [3576] = 8'd140;
   assign soundFileAmplitudes [3577] = 8'd113;
   assign soundFileAmplitudes [3578] = 8'd132;
   assign soundFileAmplitudes [3579] = 8'd141;
   assign soundFileAmplitudes [3580] = 8'd151;
   assign soundFileAmplitudes [3581] = 8'd169;
   assign soundFileAmplitudes [3582] = 8'd156;
   assign soundFileAmplitudes [3583] = 8'd130;
   assign soundFileAmplitudes [3584] = 8'd139;
   assign soundFileAmplitudes [3585] = 8'd148;
   assign soundFileAmplitudes [3586] = 8'd122;
   assign soundFileAmplitudes [3587] = 8'd117;
   assign soundFileAmplitudes [3588] = 8'd111;
   assign soundFileAmplitudes [3589] = 8'd113;
   assign soundFileAmplitudes [3590] = 8'd110;
   assign soundFileAmplitudes [3591] = 8'd93;
   assign soundFileAmplitudes [3592] = 8'd94;
   assign soundFileAmplitudes [3593] = 8'd107;
   assign soundFileAmplitudes [3594] = 8'd117;
   assign soundFileAmplitudes [3595] = 8'd108;
   assign soundFileAmplitudes [3596] = 8'd112;
   assign soundFileAmplitudes [3597] = 8'd125;
   assign soundFileAmplitudes [3598] = 8'd131;
   assign soundFileAmplitudes [3599] = 8'd134;
   assign soundFileAmplitudes [3600] = 8'd120;
   assign soundFileAmplitudes [3601] = 8'd125;
   assign soundFileAmplitudes [3602] = 8'd127;
   assign soundFileAmplitudes [3603] = 8'd133;
   assign soundFileAmplitudes [3604] = 8'd139;
   assign soundFileAmplitudes [3605] = 8'd135;
   assign soundFileAmplitudes [3606] = 8'd138;
   assign soundFileAmplitudes [3607] = 8'd136;
   assign soundFileAmplitudes [3608] = 8'd138;
   assign soundFileAmplitudes [3609] = 8'd149;
   assign soundFileAmplitudes [3610] = 8'd158;
   assign soundFileAmplitudes [3611] = 8'd157;
   assign soundFileAmplitudes [3612] = 8'd146;
   assign soundFileAmplitudes [3613] = 8'd137;
   assign soundFileAmplitudes [3614] = 8'd128;
   assign soundFileAmplitudes [3615] = 8'd123;
   assign soundFileAmplitudes [3616] = 8'd128;
   assign soundFileAmplitudes [3617] = 8'd115;
   assign soundFileAmplitudes [3618] = 8'd107;
   assign soundFileAmplitudes [3619] = 8'd114;
   assign soundFileAmplitudes [3620] = 8'd127;
   assign soundFileAmplitudes [3621] = 8'd136;
   assign soundFileAmplitudes [3622] = 8'd131;
   assign soundFileAmplitudes [3623] = 8'd122;
   assign soundFileAmplitudes [3624] = 8'd118;
   assign soundFileAmplitudes [3625] = 8'd106;
   assign soundFileAmplitudes [3626] = 8'd97;
   assign soundFileAmplitudes [3627] = 8'd113;
   assign soundFileAmplitudes [3628] = 8'd127;
   assign soundFileAmplitudes [3629] = 8'd120;
   assign soundFileAmplitudes [3630] = 8'd112;
   assign soundFileAmplitudes [3631] = 8'd87;
   assign soundFileAmplitudes [3632] = 8'd60;
   assign soundFileAmplitudes [3633] = 8'd80;
   assign soundFileAmplitudes [3634] = 8'd94;
   assign soundFileAmplitudes [3635] = 8'd105;
   assign soundFileAmplitudes [3636] = 8'd115;
   assign soundFileAmplitudes [3637] = 8'd118;
   assign soundFileAmplitudes [3638] = 8'd136;
   assign soundFileAmplitudes [3639] = 8'd155;
   assign soundFileAmplitudes [3640] = 8'd160;
   assign soundFileAmplitudes [3641] = 8'd156;
   assign soundFileAmplitudes [3642] = 8'd161;
   assign soundFileAmplitudes [3643] = 8'd166;
   assign soundFileAmplitudes [3644] = 8'd172;
   assign soundFileAmplitudes [3645] = 8'd161;
   assign soundFileAmplitudes [3646] = 8'd144;
   assign soundFileAmplitudes [3647] = 8'd134;
   assign soundFileAmplitudes [3648] = 8'd118;
   assign soundFileAmplitudes [3649] = 8'd108;
   assign soundFileAmplitudes [3650] = 8'd112;
   assign soundFileAmplitudes [3651] = 8'd128;
   assign soundFileAmplitudes [3652] = 8'd139;
   assign soundFileAmplitudes [3653] = 8'd119;
   assign soundFileAmplitudes [3654] = 8'd106;
   assign soundFileAmplitudes [3655] = 8'd120;
   assign soundFileAmplitudes [3656] = 8'd138;
   assign soundFileAmplitudes [3657] = 8'd136;
   assign soundFileAmplitudes [3658] = 8'd133;
   assign soundFileAmplitudes [3659] = 8'd141;
   assign soundFileAmplitudes [3660] = 8'd126;
   assign soundFileAmplitudes [3661] = 8'd128;
   assign soundFileAmplitudes [3662] = 8'd104;
   assign soundFileAmplitudes [3663] = 8'd76;
   assign soundFileAmplitudes [3664] = 8'd82;
   assign soundFileAmplitudes [3665] = 8'd88;
   assign soundFileAmplitudes [3666] = 8'd97;
   assign soundFileAmplitudes [3667] = 8'd106;
   assign soundFileAmplitudes [3668] = 8'd100;
   assign soundFileAmplitudes [3669] = 8'd93;
   assign soundFileAmplitudes [3670] = 8'd107;
   assign soundFileAmplitudes [3671] = 8'd115;
   assign soundFileAmplitudes [3672] = 8'd139;
   assign soundFileAmplitudes [3673] = 8'd157;
   assign soundFileAmplitudes [3674] = 8'd160;
   assign soundFileAmplitudes [3675] = 8'd177;
   assign soundFileAmplitudes [3676] = 8'd186;
   assign soundFileAmplitudes [3677] = 8'd166;
   assign soundFileAmplitudes [3678] = 8'd153;
   assign soundFileAmplitudes [3679] = 8'd143;
   assign soundFileAmplitudes [3680] = 8'd138;
   assign soundFileAmplitudes [3681] = 8'd125;
   assign soundFileAmplitudes [3682] = 8'd117;
   assign soundFileAmplitudes [3683] = 8'd123;
   assign soundFileAmplitudes [3684] = 8'd119;
   assign soundFileAmplitudes [3685] = 8'd112;
   assign soundFileAmplitudes [3686] = 8'd100;
   assign soundFileAmplitudes [3687] = 8'd106;
   assign soundFileAmplitudes [3688] = 8'd125;
   assign soundFileAmplitudes [3689] = 8'd137;
   assign soundFileAmplitudes [3690] = 8'd126;
   assign soundFileAmplitudes [3691] = 8'd130;
   assign soundFileAmplitudes [3692] = 8'd143;
   assign soundFileAmplitudes [3693] = 8'd156;
   assign soundFileAmplitudes [3694] = 8'd140;
   assign soundFileAmplitudes [3695] = 8'd118;
   assign soundFileAmplitudes [3696] = 8'd111;
   assign soundFileAmplitudes [3697] = 8'd105;
   assign soundFileAmplitudes [3698] = 8'd105;
   assign soundFileAmplitudes [3699] = 8'd93;
   assign soundFileAmplitudes [3700] = 8'd88;
   assign soundFileAmplitudes [3701] = 8'd101;
   assign soundFileAmplitudes [3702] = 8'd108;
   assign soundFileAmplitudes [3703] = 8'd107;
   assign soundFileAmplitudes [3704] = 8'd111;
   assign soundFileAmplitudes [3705] = 8'd119;
   assign soundFileAmplitudes [3706] = 8'd127;
   assign soundFileAmplitudes [3707] = 8'd131;
   assign soundFileAmplitudes [3708] = 8'd149;
   assign soundFileAmplitudes [3709] = 8'd146;
   assign soundFileAmplitudes [3710] = 8'd145;
   assign soundFileAmplitudes [3711] = 8'd151;
   assign soundFileAmplitudes [3712] = 8'd157;
   assign soundFileAmplitudes [3713] = 8'd161;
   assign soundFileAmplitudes [3714] = 8'd166;
   assign soundFileAmplitudes [3715] = 8'd166;
   assign soundFileAmplitudes [3716] = 8'd151;
   assign soundFileAmplitudes [3717] = 8'd133;
   assign soundFileAmplitudes [3718] = 8'd114;
   assign soundFileAmplitudes [3719] = 8'd107;
   assign soundFileAmplitudes [3720] = 8'd116;
   assign soundFileAmplitudes [3721] = 8'd122;
   assign soundFileAmplitudes [3722] = 8'd106;
   assign soundFileAmplitudes [3723] = 8'd121;
   assign soundFileAmplitudes [3724] = 8'd132;
   assign soundFileAmplitudes [3725] = 8'd138;
   assign soundFileAmplitudes [3726] = 8'd138;
   assign soundFileAmplitudes [3727] = 8'd97;
   assign soundFileAmplitudes [3728] = 8'd81;
   assign soundFileAmplitudes [3729] = 8'd93;
   assign soundFileAmplitudes [3730] = 8'd108;
   assign soundFileAmplitudes [3731] = 8'd120;
   assign soundFileAmplitudes [3732] = 8'd113;
   assign soundFileAmplitudes [3733] = 8'd110;
   assign soundFileAmplitudes [3734] = 8'd113;
   assign soundFileAmplitudes [3735] = 8'd121;
   assign soundFileAmplitudes [3736] = 8'd119;
   assign soundFileAmplitudes [3737] = 8'd124;
   assign soundFileAmplitudes [3738] = 8'd145;
   assign soundFileAmplitudes [3739] = 8'd145;
   assign soundFileAmplitudes [3740] = 8'd134;
   assign soundFileAmplitudes [3741] = 8'd134;
   assign soundFileAmplitudes [3742] = 8'd130;
   assign soundFileAmplitudes [3743] = 8'd122;
   assign soundFileAmplitudes [3744] = 8'd133;
   assign soundFileAmplitudes [3745] = 8'd139;
   assign soundFileAmplitudes [3746] = 8'd142;
   assign soundFileAmplitudes [3747] = 8'd151;
   assign soundFileAmplitudes [3748] = 8'd149;
   assign soundFileAmplitudes [3749] = 8'd133;
   assign soundFileAmplitudes [3750] = 8'd133;
   assign soundFileAmplitudes [3751] = 8'd140;
   assign soundFileAmplitudes [3752] = 8'd145;
   assign soundFileAmplitudes [3753] = 8'd138;
   assign soundFileAmplitudes [3754] = 8'd123;
   assign soundFileAmplitudes [3755] = 8'd115;
   assign soundFileAmplitudes [3756] = 8'd95;
   assign soundFileAmplitudes [3757] = 8'd105;
   assign soundFileAmplitudes [3758] = 8'd105;
   assign soundFileAmplitudes [3759] = 8'd91;
   assign soundFileAmplitudes [3760] = 8'd90;
   assign soundFileAmplitudes [3761] = 8'd86;
   assign soundFileAmplitudes [3762] = 8'd86;
   assign soundFileAmplitudes [3763] = 8'd104;
   assign soundFileAmplitudes [3764] = 8'd115;
   assign soundFileAmplitudes [3765] = 8'd117;
   assign soundFileAmplitudes [3766] = 8'd134;
   assign soundFileAmplitudes [3767] = 8'd139;
   assign soundFileAmplitudes [3768] = 8'd145;
   assign soundFileAmplitudes [3769] = 8'd135;
   assign soundFileAmplitudes [3770] = 8'd163;
   assign soundFileAmplitudes [3771] = 8'd166;
   assign soundFileAmplitudes [3772] = 8'd158;
   assign soundFileAmplitudes [3773] = 8'd149;
   assign soundFileAmplitudes [3774] = 8'd129;
   assign soundFileAmplitudes [3775] = 8'd142;
   assign soundFileAmplitudes [3776] = 8'd132;
   assign soundFileAmplitudes [3777] = 8'd130;
   assign soundFileAmplitudes [3778] = 8'd135;
   assign soundFileAmplitudes [3779] = 8'd129;
   assign soundFileAmplitudes [3780] = 8'd110;
   assign soundFileAmplitudes [3781] = 8'd110;
   assign soundFileAmplitudes [3782] = 8'd114;
   assign soundFileAmplitudes [3783] = 8'd117;
   assign soundFileAmplitudes [3784] = 8'd117;
   assign soundFileAmplitudes [3785] = 8'd119;
   assign soundFileAmplitudes [3786] = 8'd113;
   assign soundFileAmplitudes [3787] = 8'd123;
   assign soundFileAmplitudes [3788] = 8'd142;
   assign soundFileAmplitudes [3789] = 8'd133;
   assign soundFileAmplitudes [3790] = 8'd141;
   assign soundFileAmplitudes [3791] = 8'd135;
   assign soundFileAmplitudes [3792] = 8'd99;
   assign soundFileAmplitudes [3793] = 8'd80;
   assign soundFileAmplitudes [3794] = 8'd72;
   assign soundFileAmplitudes [3795] = 8'd78;
   assign soundFileAmplitudes [3796] = 8'd103;
   assign soundFileAmplitudes [3797] = 8'd111;
   assign soundFileAmplitudes [3798] = 8'd116;
   assign soundFileAmplitudes [3799] = 8'd115;
   assign soundFileAmplitudes [3800] = 8'd116;
   assign soundFileAmplitudes [3801] = 8'd139;
   assign soundFileAmplitudes [3802] = 8'd174;
   assign soundFileAmplitudes [3803] = 8'd186;
   assign soundFileAmplitudes [3804] = 8'd192;
   assign soundFileAmplitudes [3805] = 8'd175;
   assign soundFileAmplitudes [3806] = 8'd160;
   assign soundFileAmplitudes [3807] = 8'd147;
   assign soundFileAmplitudes [3808] = 8'd145;
   assign soundFileAmplitudes [3809] = 8'd157;
   assign soundFileAmplitudes [3810] = 8'd138;
   assign soundFileAmplitudes [3811] = 8'd134;
   assign soundFileAmplitudes [3812] = 8'd109;
   assign soundFileAmplitudes [3813] = 8'd91;
   assign soundFileAmplitudes [3814] = 8'd82;
   assign soundFileAmplitudes [3815] = 8'd72;
   assign soundFileAmplitudes [3816] = 8'd80;
   assign soundFileAmplitudes [3817] = 8'd89;
   assign soundFileAmplitudes [3818] = 8'd91;
   assign soundFileAmplitudes [3819] = 8'd106;
   assign soundFileAmplitudes [3820] = 8'd133;
   assign soundFileAmplitudes [3821] = 8'd151;
   assign soundFileAmplitudes [3822] = 8'd159;
   assign soundFileAmplitudes [3823] = 8'd143;
   assign soundFileAmplitudes [3824] = 8'd107;
   assign soundFileAmplitudes [3825] = 8'd106;
   assign soundFileAmplitudes [3826] = 8'd118;
   assign soundFileAmplitudes [3827] = 8'd121;
   assign soundFileAmplitudes [3828] = 8'd124;
   assign soundFileAmplitudes [3829] = 8'd110;
   assign soundFileAmplitudes [3830] = 8'd97;
   assign soundFileAmplitudes [3831] = 8'd92;
   assign soundFileAmplitudes [3832] = 8'd104;
   assign soundFileAmplitudes [3833] = 8'd130;
   assign soundFileAmplitudes [3834] = 8'd152;
   assign soundFileAmplitudes [3835] = 8'd165;
   assign soundFileAmplitudes [3836] = 8'd168;
   assign soundFileAmplitudes [3837] = 8'd163;
   assign soundFileAmplitudes [3838] = 8'd170;
   assign soundFileAmplitudes [3839] = 8'd177;
   assign soundFileAmplitudes [3840] = 8'd194;
   assign soundFileAmplitudes [3841] = 8'd190;
   assign soundFileAmplitudes [3842] = 8'd152;
   assign soundFileAmplitudes [3843] = 8'd144;
   assign soundFileAmplitudes [3844] = 8'd143;
   assign soundFileAmplitudes [3845] = 8'd118;
   assign soundFileAmplitudes [3846] = 8'd116;
   assign soundFileAmplitudes [3847] = 8'd111;
   assign soundFileAmplitudes [3848] = 8'd91;
   assign soundFileAmplitudes [3849] = 8'd85;
   assign soundFileAmplitudes [3850] = 8'd75;
   assign soundFileAmplitudes [3851] = 8'd85;
   assign soundFileAmplitudes [3852] = 8'd81;
   assign soundFileAmplitudes [3853] = 8'd83;
   assign soundFileAmplitudes [3854] = 8'd90;
   assign soundFileAmplitudes [3855] = 8'd100;
   assign soundFileAmplitudes [3856] = 8'd111;
   assign soundFileAmplitudes [3857] = 8'd98;
   assign soundFileAmplitudes [3858] = 8'd99;
   assign soundFileAmplitudes [3859] = 8'd102;
   assign soundFileAmplitudes [3860] = 8'd112;
   assign soundFileAmplitudes [3861] = 8'd119;
   assign soundFileAmplitudes [3862] = 8'd119;
   assign soundFileAmplitudes [3863] = 8'd134;
   assign soundFileAmplitudes [3864] = 8'd140;
   assign soundFileAmplitudes [3865] = 8'd137;
   assign soundFileAmplitudes [3866] = 8'd140;
   assign soundFileAmplitudes [3867] = 8'd150;
   assign soundFileAmplitudes [3868] = 8'd161;
   assign soundFileAmplitudes [3869] = 8'd165;
   assign soundFileAmplitudes [3870] = 8'd155;
   assign soundFileAmplitudes [3871] = 8'd149;
   assign soundFileAmplitudes [3872] = 8'd155;
   assign soundFileAmplitudes [3873] = 8'd156;
   assign soundFileAmplitudes [3874] = 8'd164;
   assign soundFileAmplitudes [3875] = 8'd154;
   assign soundFileAmplitudes [3876] = 8'd161;
   assign soundFileAmplitudes [3877] = 8'd163;
   assign soundFileAmplitudes [3878] = 8'd152;
   assign soundFileAmplitudes [3879] = 8'd138;
   assign soundFileAmplitudes [3880] = 8'd114;
   assign soundFileAmplitudes [3881] = 8'd104;
   assign soundFileAmplitudes [3882] = 8'd103;
   assign soundFileAmplitudes [3883] = 8'd98;
   assign soundFileAmplitudes [3884] = 8'd87;
   assign soundFileAmplitudes [3885] = 8'd109;
   assign soundFileAmplitudes [3886] = 8'd124;
   assign soundFileAmplitudes [3887] = 8'd133;
   assign soundFileAmplitudes [3888] = 8'd111;
   assign soundFileAmplitudes [3889] = 8'd91;
   assign soundFileAmplitudes [3890] = 8'd75;
   assign soundFileAmplitudes [3891] = 8'd64;
   assign soundFileAmplitudes [3892] = 8'd75;
   assign soundFileAmplitudes [3893] = 8'd84;
   assign soundFileAmplitudes [3894] = 8'd98;
   assign soundFileAmplitudes [3895] = 8'd111;
   assign soundFileAmplitudes [3896] = 8'd132;
   assign soundFileAmplitudes [3897] = 8'd134;
   assign soundFileAmplitudes [3898] = 8'd129;
   assign soundFileAmplitudes [3899] = 8'd127;
   assign soundFileAmplitudes [3900] = 8'd143;
   assign soundFileAmplitudes [3901] = 8'd168;
   assign soundFileAmplitudes [3902] = 8'd164;
   assign soundFileAmplitudes [3903] = 8'd159;
   assign soundFileAmplitudes [3904] = 8'd156;
   assign soundFileAmplitudes [3905] = 8'd154;
   assign soundFileAmplitudes [3906] = 8'd156;
   assign soundFileAmplitudes [3907] = 8'd148;
   assign soundFileAmplitudes [3908] = 8'd147;
   assign soundFileAmplitudes [3909] = 8'd153;
   assign soundFileAmplitudes [3910] = 8'd161;
   assign soundFileAmplitudes [3911] = 8'd151;
   assign soundFileAmplitudes [3912] = 8'd139;
   assign soundFileAmplitudes [3913] = 8'd106;
   assign soundFileAmplitudes [3914] = 8'd87;
   assign soundFileAmplitudes [3915] = 8'd110;
   assign soundFileAmplitudes [3916] = 8'd110;
   assign soundFileAmplitudes [3917] = 8'd103;
   assign soundFileAmplitudes [3918] = 8'd99;
   assign soundFileAmplitudes [3919] = 8'd109;
   assign soundFileAmplitudes [3920] = 8'd115;
   assign soundFileAmplitudes [3921] = 8'd127;
   assign soundFileAmplitudes [3922] = 8'd101;
   assign soundFileAmplitudes [3923] = 8'd66;
   assign soundFileAmplitudes [3924] = 8'd81;
   assign soundFileAmplitudes [3925] = 8'd109;
   assign soundFileAmplitudes [3926] = 8'd143;
   assign soundFileAmplitudes [3927] = 8'd120;
   assign soundFileAmplitudes [3928] = 8'd96;
   assign soundFileAmplitudes [3929] = 8'd103;
   assign soundFileAmplitudes [3930] = 8'd101;
   assign soundFileAmplitudes [3931] = 8'd115;
   assign soundFileAmplitudes [3932] = 8'd116;
   assign soundFileAmplitudes [3933] = 8'd135;
   assign soundFileAmplitudes [3934] = 8'd157;
   assign soundFileAmplitudes [3935] = 8'd168;
   assign soundFileAmplitudes [3936] = 8'd163;
   assign soundFileAmplitudes [3937] = 8'd138;
   assign soundFileAmplitudes [3938] = 8'd126;
   assign soundFileAmplitudes [3939] = 8'd124;
   assign soundFileAmplitudes [3940] = 8'd134;
   assign soundFileAmplitudes [3941] = 8'd147;
   assign soundFileAmplitudes [3942] = 8'd149;
   assign soundFileAmplitudes [3943] = 8'd167;
   assign soundFileAmplitudes [3944] = 8'd152;
   assign soundFileAmplitudes [3945] = 8'd137;
   assign soundFileAmplitudes [3946] = 8'd136;
   assign soundFileAmplitudes [3947] = 8'd136;
   assign soundFileAmplitudes [3948] = 8'd146;
   assign soundFileAmplitudes [3949] = 8'd135;
   assign soundFileAmplitudes [3950] = 8'd120;
   assign soundFileAmplitudes [3951] = 8'd114;
   assign soundFileAmplitudes [3952] = 8'd117;
   assign soundFileAmplitudes [3953] = 8'd120;
   assign soundFileAmplitudes [3954] = 8'd133;
   assign soundFileAmplitudes [3955] = 8'd109;
   assign soundFileAmplitudes [3956] = 8'd91;
   assign soundFileAmplitudes [3957] = 8'd81;
   assign soundFileAmplitudes [3958] = 8'd95;
   assign soundFileAmplitudes [3959] = 8'd119;
   assign soundFileAmplitudes [3960] = 8'd128;
   assign soundFileAmplitudes [3961] = 8'd117;
   assign soundFileAmplitudes [3962] = 8'd123;
   assign soundFileAmplitudes [3963] = 8'd141;
   assign soundFileAmplitudes [3964] = 8'd144;
   assign soundFileAmplitudes [3965] = 8'd158;
   assign soundFileAmplitudes [3966] = 8'd136;
   assign soundFileAmplitudes [3967] = 8'd136;
   assign soundFileAmplitudes [3968] = 8'd131;
   assign soundFileAmplitudes [3969] = 8'd129;
   assign soundFileAmplitudes [3970] = 8'd126;
   assign soundFileAmplitudes [3971] = 8'd120;
   assign soundFileAmplitudes [3972] = 8'd117;
   assign soundFileAmplitudes [3973] = 8'd113;
   assign soundFileAmplitudes [3974] = 8'd111;
   assign soundFileAmplitudes [3975] = 8'd111;
   assign soundFileAmplitudes [3976] = 8'd111;
   assign soundFileAmplitudes [3977] = 8'd105;
   assign soundFileAmplitudes [3978] = 8'd114;
   assign soundFileAmplitudes [3979] = 8'd108;
   assign soundFileAmplitudes [3980] = 8'd115;
   assign soundFileAmplitudes [3981] = 8'd140;
   assign soundFileAmplitudes [3982] = 8'd154;
   assign soundFileAmplitudes [3983] = 8'd143;
   assign soundFileAmplitudes [3984] = 8'd140;
   assign soundFileAmplitudes [3985] = 8'd113;
   assign soundFileAmplitudes [3986] = 8'd124;
   assign soundFileAmplitudes [3987] = 8'd135;
   assign soundFileAmplitudes [3988] = 8'd107;
   assign soundFileAmplitudes [3989] = 8'd100;
   assign soundFileAmplitudes [3990] = 8'd106;
   assign soundFileAmplitudes [3991] = 8'd123;
   assign soundFileAmplitudes [3992] = 8'd130;
   assign soundFileAmplitudes [3993] = 8'd137;
   assign soundFileAmplitudes [3994] = 8'd143;
   assign soundFileAmplitudes [3995] = 8'd137;
   assign soundFileAmplitudes [3996] = 8'd140;
   assign soundFileAmplitudes [3997] = 8'd161;
   assign soundFileAmplitudes [3998] = 8'd177;
   assign soundFileAmplitudes [3999] = 8'd185;
   assign soundFileAmplitudes [4000] = 8'd167;
   assign soundFileAmplitudes [4001] = 8'd166;
   assign soundFileAmplitudes [4002] = 8'd167;
   assign soundFileAmplitudes [4003] = 8'd171;
   assign soundFileAmplitudes [4004] = 8'd148;
   assign soundFileAmplitudes [4005] = 8'd103;
   assign soundFileAmplitudes [4006] = 8'd95;
   assign soundFileAmplitudes [4007] = 8'd82;
   assign soundFileAmplitudes [4008] = 8'd80;
   assign soundFileAmplitudes [4009] = 8'd72;
   assign soundFileAmplitudes [4010] = 8'd61;
   assign soundFileAmplitudes [4011] = 8'd67;
   assign soundFileAmplitudes [4012] = 8'd84;
   assign soundFileAmplitudes [4013] = 8'd103;
   assign soundFileAmplitudes [4014] = 8'd111;
   assign soundFileAmplitudes [4015] = 8'd99;
   assign soundFileAmplitudes [4016] = 8'd93;
   assign soundFileAmplitudes [4017] = 8'd120;
   assign soundFileAmplitudes [4018] = 8'd130;
   assign soundFileAmplitudes [4019] = 8'd143;
   assign soundFileAmplitudes [4020] = 8'd124;
   assign soundFileAmplitudes [4021] = 8'd83;
   assign soundFileAmplitudes [4022] = 8'd101;
   assign soundFileAmplitudes [4023] = 8'd105;
   assign soundFileAmplitudes [4024] = 8'd116;
   assign soundFileAmplitudes [4025] = 8'd144;
   assign soundFileAmplitudes [4026] = 8'd149;
   assign soundFileAmplitudes [4027] = 8'd147;
   assign soundFileAmplitudes [4028] = 8'd152;
   assign soundFileAmplitudes [4029] = 8'd163;
   assign soundFileAmplitudes [4030] = 8'd170;
   assign soundFileAmplitudes [4031] = 8'd178;
   assign soundFileAmplitudes [4032] = 8'd184;
   assign soundFileAmplitudes [4033] = 8'd176;
   assign soundFileAmplitudes [4034] = 8'd169;
   assign soundFileAmplitudes [4035] = 8'd171;
   assign soundFileAmplitudes [4036] = 8'd156;
   assign soundFileAmplitudes [4037] = 8'd142;
   assign soundFileAmplitudes [4038] = 8'd146;
   assign soundFileAmplitudes [4039] = 8'd140;
   assign soundFileAmplitudes [4040] = 8'd116;
   assign soundFileAmplitudes [4041] = 8'd128;
   assign soundFileAmplitudes [4042] = 8'd119;
   assign soundFileAmplitudes [4043] = 8'd101;
   assign soundFileAmplitudes [4044] = 8'd82;
   assign soundFileAmplitudes [4045] = 8'd40;
   assign soundFileAmplitudes [4046] = 8'd46;
   assign soundFileAmplitudes [4047] = 8'd58;
   assign soundFileAmplitudes [4048] = 8'd65;
   assign soundFileAmplitudes [4049] = 8'd86;
   assign soundFileAmplitudes [4050] = 8'd101;
   assign soundFileAmplitudes [4051] = 8'd98;
   assign soundFileAmplitudes [4052] = 8'd100;
   assign soundFileAmplitudes [4053] = 8'd105;
   assign soundFileAmplitudes [4054] = 8'd106;
   assign soundFileAmplitudes [4055] = 8'd107;
   assign soundFileAmplitudes [4056] = 8'd111;
   assign soundFileAmplitudes [4057] = 8'd140;
   assign soundFileAmplitudes [4058] = 8'd160;
   assign soundFileAmplitudes [4059] = 8'd154;
   assign soundFileAmplitudes [4060] = 8'd156;
   assign soundFileAmplitudes [4061] = 8'd154;
   assign soundFileAmplitudes [4062] = 8'd159;
   assign soundFileAmplitudes [4063] = 8'd168;
   assign soundFileAmplitudes [4064] = 8'd173;
   assign soundFileAmplitudes [4065] = 8'd166;
   assign soundFileAmplitudes [4066] = 8'd158;
   assign soundFileAmplitudes [4067] = 8'd165;
   assign soundFileAmplitudes [4068] = 8'd164;
   assign soundFileAmplitudes [4069] = 8'd165;
   assign soundFileAmplitudes [4070] = 8'd166;
   assign soundFileAmplitudes [4071] = 8'd163;
   assign soundFileAmplitudes [4072] = 8'd151;
   assign soundFileAmplitudes [4073] = 8'd140;
   assign soundFileAmplitudes [4074] = 8'd134;
   assign soundFileAmplitudes [4075] = 8'd115;
   assign soundFileAmplitudes [4076] = 8'd98;
   assign soundFileAmplitudes [4077] = 8'd88;
   assign soundFileAmplitudes [4078] = 8'd100;
   assign soundFileAmplitudes [4079] = 8'd91;
   assign soundFileAmplitudes [4080] = 8'd77;
   assign soundFileAmplitudes [4081] = 8'd71;
   assign soundFileAmplitudes [4082] = 8'd78;
   assign soundFileAmplitudes [4083] = 8'd105;
   assign soundFileAmplitudes [4084] = 8'd85;
   assign soundFileAmplitudes [4085] = 8'd71;
   assign soundFileAmplitudes [4086] = 8'd68;
   assign soundFileAmplitudes [4087] = 8'd66;
   assign soundFileAmplitudes [4088] = 8'd79;
   assign soundFileAmplitudes [4089] = 8'd112;
   assign soundFileAmplitudes [4090] = 8'd127;
   assign soundFileAmplitudes [4091] = 8'd131;
   assign soundFileAmplitudes [4092] = 8'd120;
   assign soundFileAmplitudes [4093] = 8'd122;
   assign soundFileAmplitudes [4094] = 8'd145;
   assign soundFileAmplitudes [4095] = 8'd160;
   assign soundFileAmplitudes [4096] = 8'd187;
   assign soundFileAmplitudes [4097] = 8'd187;
   assign soundFileAmplitudes [4098] = 8'd172;
   assign soundFileAmplitudes [4099] = 8'd156;
   assign soundFileAmplitudes [4100] = 8'd159;
   assign soundFileAmplitudes [4101] = 8'd165;
   assign soundFileAmplitudes [4102] = 8'd163;
   assign soundFileAmplitudes [4103] = 8'd158;
   assign soundFileAmplitudes [4104] = 8'd155;
   assign soundFileAmplitudes [4105] = 8'd157;
   assign soundFileAmplitudes [4106] = 8'd160;
   assign soundFileAmplitudes [4107] = 8'd157;
   assign soundFileAmplitudes [4108] = 8'd142;
   assign soundFileAmplitudes [4109] = 8'd123;
   assign soundFileAmplitudes [4110] = 8'd113;
   assign soundFileAmplitudes [4111] = 8'd114;
   assign soundFileAmplitudes [4112] = 8'd118;
   assign soundFileAmplitudes [4113] = 8'd105;
   assign soundFileAmplitudes [4114] = 8'd90;
   assign soundFileAmplitudes [4115] = 8'd99;
   assign soundFileAmplitudes [4116] = 8'd95;
   assign soundFileAmplitudes [4117] = 8'd99;
   assign soundFileAmplitudes [4118] = 8'd79;
   assign soundFileAmplitudes [4119] = 8'd50;
   assign soundFileAmplitudes [4120] = 8'd61;
   assign soundFileAmplitudes [4121] = 8'd83;
   assign soundFileAmplitudes [4122] = 8'd120;
   assign soundFileAmplitudes [4123] = 8'd138;
   assign soundFileAmplitudes [4124] = 8'd118;
   assign soundFileAmplitudes [4125] = 8'd113;
   assign soundFileAmplitudes [4126] = 8'd130;
   assign soundFileAmplitudes [4127] = 8'd144;
   assign soundFileAmplitudes [4128] = 8'd144;
   assign soundFileAmplitudes [4129] = 8'd133;
   assign soundFileAmplitudes [4130] = 8'd127;
   assign soundFileAmplitudes [4131] = 8'd126;
   assign soundFileAmplitudes [4132] = 8'd139;
   assign soundFileAmplitudes [4133] = 8'd158;
   assign soundFileAmplitudes [4134] = 8'd164;
   assign soundFileAmplitudes [4135] = 8'd158;
   assign soundFileAmplitudes [4136] = 8'd162;
   assign soundFileAmplitudes [4137] = 8'd155;
   assign soundFileAmplitudes [4138] = 8'd157;
   assign soundFileAmplitudes [4139] = 8'd169;
   assign soundFileAmplitudes [4140] = 8'd164;
   assign soundFileAmplitudes [4141] = 8'd147;
   assign soundFileAmplitudes [4142] = 8'd130;
   assign soundFileAmplitudes [4143] = 8'd125;
   assign soundFileAmplitudes [4144] = 8'd116;
   assign soundFileAmplitudes [4145] = 8'd110;
   assign soundFileAmplitudes [4146] = 8'd108;
   assign soundFileAmplitudes [4147] = 8'd113;
   assign soundFileAmplitudes [4148] = 8'd117;
   assign soundFileAmplitudes [4149] = 8'd119;
   assign soundFileAmplitudes [4150] = 8'd115;
   assign soundFileAmplitudes [4151] = 8'd93;
   assign soundFileAmplitudes [4152] = 8'd72;
   assign soundFileAmplitudes [4153] = 8'd57;
   assign soundFileAmplitudes [4154] = 8'd52;
   assign soundFileAmplitudes [4155] = 8'd86;
   assign soundFileAmplitudes [4156] = 8'd128;
   assign soundFileAmplitudes [4157] = 8'd143;
   assign soundFileAmplitudes [4158] = 8'd125;
   assign soundFileAmplitudes [4159] = 8'd124;
   assign soundFileAmplitudes [4160] = 8'd129;
   assign soundFileAmplitudes [4161] = 8'd161;
   assign soundFileAmplitudes [4162] = 8'd187;
   assign soundFileAmplitudes [4163] = 8'd154;
   assign soundFileAmplitudes [4164] = 8'd135;
   assign soundFileAmplitudes [4165] = 8'd114;
   assign soundFileAmplitudes [4166] = 8'd121;
   assign soundFileAmplitudes [4167] = 8'd122;
   assign soundFileAmplitudes [4168] = 8'd111;
   assign soundFileAmplitudes [4169] = 8'd115;
   assign soundFileAmplitudes [4170] = 8'd126;
   assign soundFileAmplitudes [4171] = 8'd145;
   assign soundFileAmplitudes [4172] = 8'd151;
   assign soundFileAmplitudes [4173] = 8'd134;
   assign soundFileAmplitudes [4174] = 8'd130;
   assign soundFileAmplitudes [4175] = 8'd129;
   assign soundFileAmplitudes [4176] = 8'd124;
   assign soundFileAmplitudes [4177] = 8'd138;
   assign soundFileAmplitudes [4178] = 8'd140;
   assign soundFileAmplitudes [4179] = 8'd140;
   assign soundFileAmplitudes [4180] = 8'd140;
   assign soundFileAmplitudes [4181] = 8'd136;
   assign soundFileAmplitudes [4182] = 8'd126;
   assign soundFileAmplitudes [4183] = 8'd135;
   assign soundFileAmplitudes [4184] = 8'd129;
   assign soundFileAmplitudes [4185] = 8'd112;
   assign soundFileAmplitudes [4186] = 8'd108;
   assign soundFileAmplitudes [4187] = 8'd103;
   assign soundFileAmplitudes [4188] = 8'd101;
   assign soundFileAmplitudes [4189] = 8'd104;
   assign soundFileAmplitudes [4190] = 8'd91;
   assign soundFileAmplitudes [4191] = 8'd84;
   assign soundFileAmplitudes [4192] = 8'd97;
   assign soundFileAmplitudes [4193] = 8'd114;
   assign soundFileAmplitudes [4194] = 8'd137;
   assign soundFileAmplitudes [4195] = 8'd146;
   assign soundFileAmplitudes [4196] = 8'd138;
   assign soundFileAmplitudes [4197] = 8'd127;
   assign soundFileAmplitudes [4198] = 8'd155;
   assign soundFileAmplitudes [4199] = 8'd167;
   assign soundFileAmplitudes [4200] = 8'd175;
   assign soundFileAmplitudes [4201] = 8'd138;
   assign soundFileAmplitudes [4202] = 8'd98;
   assign soundFileAmplitudes [4203] = 8'd114;
   assign soundFileAmplitudes [4204] = 8'd115;
   assign soundFileAmplitudes [4205] = 8'd125;
   assign soundFileAmplitudes [4206] = 8'd116;
   assign soundFileAmplitudes [4207] = 8'd100;
   assign soundFileAmplitudes [4208] = 8'd101;
   assign soundFileAmplitudes [4209] = 8'd106;
   assign soundFileAmplitudes [4210] = 8'd120;
   assign soundFileAmplitudes [4211] = 8'd136;
   assign soundFileAmplitudes [4212] = 8'd125;
   assign soundFileAmplitudes [4213] = 8'd130;
   assign soundFileAmplitudes [4214] = 8'd155;
   assign soundFileAmplitudes [4215] = 8'd149;
   assign soundFileAmplitudes [4216] = 8'd150;
   assign soundFileAmplitudes [4217] = 8'd144;
   assign soundFileAmplitudes [4218] = 8'd129;
   assign soundFileAmplitudes [4219] = 8'd121;
   assign soundFileAmplitudes [4220] = 8'd107;
   assign soundFileAmplitudes [4221] = 8'd109;
   assign soundFileAmplitudes [4222] = 8'd128;
   assign soundFileAmplitudes [4223] = 8'd138;
   assign soundFileAmplitudes [4224] = 8'd134;
   assign soundFileAmplitudes [4225] = 8'd123;
   assign soundFileAmplitudes [4226] = 8'd110;
   assign soundFileAmplitudes [4227] = 8'd90;
   assign soundFileAmplitudes [4228] = 8'd90;
   assign soundFileAmplitudes [4229] = 8'd113;
   assign soundFileAmplitudes [4230] = 8'd129;
   assign soundFileAmplitudes [4231] = 8'd136;
   assign soundFileAmplitudes [4232] = 8'd138;
   assign soundFileAmplitudes [4233] = 8'd151;
   assign soundFileAmplitudes [4234] = 8'd144;
   assign soundFileAmplitudes [4235] = 8'd136;
   assign soundFileAmplitudes [4236] = 8'd146;
   assign soundFileAmplitudes [4237] = 8'd151;
   assign soundFileAmplitudes [4238] = 8'd146;
   assign soundFileAmplitudes [4239] = 8'd127;
   assign soundFileAmplitudes [4240] = 8'd106;
   assign soundFileAmplitudes [4241] = 8'd107;
   assign soundFileAmplitudes [4242] = 8'd110;
   assign soundFileAmplitudes [4243] = 8'd96;
   assign soundFileAmplitudes [4244] = 8'd94;
   assign soundFileAmplitudes [4245] = 8'd98;
   assign soundFileAmplitudes [4246] = 8'd111;
   assign soundFileAmplitudes [4247] = 8'd129;
   assign soundFileAmplitudes [4248] = 8'd139;
   assign soundFileAmplitudes [4249] = 8'd144;
   assign soundFileAmplitudes [4250] = 8'd146;
   assign soundFileAmplitudes [4251] = 8'd149;
   assign soundFileAmplitudes [4252] = 8'd142;
   assign soundFileAmplitudes [4253] = 8'd133;
   assign soundFileAmplitudes [4254] = 8'd124;
   assign soundFileAmplitudes [4255] = 8'd124;
   assign soundFileAmplitudes [4256] = 8'd135;
   assign soundFileAmplitudes [4257] = 8'd131;
   assign soundFileAmplitudes [4258] = 8'd131;
   assign soundFileAmplitudes [4259] = 8'd131;
   assign soundFileAmplitudes [4260] = 8'd129;
   assign soundFileAmplitudes [4261] = 8'd120;
   assign soundFileAmplitudes [4262] = 8'd118;
   assign soundFileAmplitudes [4263] = 8'd109;
   assign soundFileAmplitudes [4264] = 8'd105;
   assign soundFileAmplitudes [4265] = 8'd122;
   assign soundFileAmplitudes [4266] = 8'd125;
   assign soundFileAmplitudes [4267] = 8'd136;
   assign soundFileAmplitudes [4268] = 8'd131;
   assign soundFileAmplitudes [4269] = 8'd129;
   assign soundFileAmplitudes [4270] = 8'd153;
   assign soundFileAmplitudes [4271] = 8'd172;
   assign soundFileAmplitudes [4272] = 8'd170;
   assign soundFileAmplitudes [4273] = 8'd147;
   assign soundFileAmplitudes [4274] = 8'd125;
   assign soundFileAmplitudes [4275] = 8'd120;
   assign soundFileAmplitudes [4276] = 8'd131;
   assign soundFileAmplitudes [4277] = 8'd120;
   assign soundFileAmplitudes [4278] = 8'd91;
   assign soundFileAmplitudes [4279] = 8'd97;
   assign soundFileAmplitudes [4280] = 8'd103;
   assign soundFileAmplitudes [4281] = 8'd96;
   assign soundFileAmplitudes [4282] = 8'd102;
   assign soundFileAmplitudes [4283] = 8'd101;
   assign soundFileAmplitudes [4284] = 8'd103;
   assign soundFileAmplitudes [4285] = 8'd99;
   assign soundFileAmplitudes [4286] = 8'd110;
   assign soundFileAmplitudes [4287] = 8'd129;
   assign soundFileAmplitudes [4288] = 8'd135;
   assign soundFileAmplitudes [4289] = 8'd139;
   assign soundFileAmplitudes [4290] = 8'd144;
   assign soundFileAmplitudes [4291] = 8'd134;
   assign soundFileAmplitudes [4292] = 8'd125;
   assign soundFileAmplitudes [4293] = 8'd125;
   assign soundFileAmplitudes [4294] = 8'd124;
   assign soundFileAmplitudes [4295] = 8'd133;
   assign soundFileAmplitudes [4296] = 8'd125;
   assign soundFileAmplitudes [4297] = 8'd120;
   assign soundFileAmplitudes [4298] = 8'd120;
   assign soundFileAmplitudes [4299] = 8'd105;
   assign soundFileAmplitudes [4300] = 8'd106;
   assign soundFileAmplitudes [4301] = 8'd119;
   assign soundFileAmplitudes [4302] = 8'd132;
   assign soundFileAmplitudes [4303] = 8'd142;
   assign soundFileAmplitudes [4304] = 8'd149;
   assign soundFileAmplitudes [4305] = 8'd154;
   assign soundFileAmplitudes [4306] = 8'd160;
   assign soundFileAmplitudes [4307] = 8'd169;
   assign soundFileAmplitudes [4308] = 8'd166;
   assign soundFileAmplitudes [4309] = 8'd161;
   assign soundFileAmplitudes [4310] = 8'd149;
   assign soundFileAmplitudes [4311] = 8'd121;
   assign soundFileAmplitudes [4312] = 8'd118;
   assign soundFileAmplitudes [4313] = 8'd108;
   assign soundFileAmplitudes [4314] = 8'd114;
   assign soundFileAmplitudes [4315] = 8'd129;
   assign soundFileAmplitudes [4316] = 8'd94;
   assign soundFileAmplitudes [4317] = 8'd70;
   assign soundFileAmplitudes [4318] = 8'd73;
   assign soundFileAmplitudes [4319] = 8'd75;
   assign soundFileAmplitudes [4320] = 8'd74;
   assign soundFileAmplitudes [4321] = 8'd77;
   assign soundFileAmplitudes [4322] = 8'd97;
   assign soundFileAmplitudes [4323] = 8'd115;
   assign soundFileAmplitudes [4324] = 8'd132;
   assign soundFileAmplitudes [4325] = 8'd147;
   assign soundFileAmplitudes [4326] = 8'd145;
   assign soundFileAmplitudes [4327] = 8'd139;
   assign soundFileAmplitudes [4328] = 8'd144;
   assign soundFileAmplitudes [4329] = 8'd152;
   assign soundFileAmplitudes [4330] = 8'd145;
   assign soundFileAmplitudes [4331] = 8'd153;
   assign soundFileAmplitudes [4332] = 8'd151;
   assign soundFileAmplitudes [4333] = 8'd142;
   assign soundFileAmplitudes [4334] = 8'd131;
   assign soundFileAmplitudes [4335] = 8'd110;
   assign soundFileAmplitudes [4336] = 8'd102;
   assign soundFileAmplitudes [4337] = 8'd113;
   assign soundFileAmplitudes [4338] = 8'd129;
   assign soundFileAmplitudes [4339] = 8'd138;
   assign soundFileAmplitudes [4340] = 8'd150;
   assign soundFileAmplitudes [4341] = 8'd147;
   assign soundFileAmplitudes [4342] = 8'd143;
   assign soundFileAmplitudes [4343] = 8'd148;
   assign soundFileAmplitudes [4344] = 8'd165;
   assign soundFileAmplitudes [4345] = 8'd158;
   assign soundFileAmplitudes [4346] = 8'd147;
   assign soundFileAmplitudes [4347] = 8'd135;
   assign soundFileAmplitudes [4348] = 8'd141;
   assign soundFileAmplitudes [4349] = 8'd125;
   assign soundFileAmplitudes [4350] = 8'd110;
   assign soundFileAmplitudes [4351] = 8'd124;
   assign soundFileAmplitudes [4352] = 8'd125;
   assign soundFileAmplitudes [4353] = 8'd133;
   assign soundFileAmplitudes [4354] = 8'd83;
   assign soundFileAmplitudes [4355] = 8'd58;
   assign soundFileAmplitudes [4356] = 8'd69;
   assign soundFileAmplitudes [4357] = 8'd71;
   assign soundFileAmplitudes [4358] = 8'd87;
   assign soundFileAmplitudes [4359] = 8'd103;
   assign soundFileAmplitudes [4360] = 8'd118;
   assign soundFileAmplitudes [4361] = 8'd125;
   assign soundFileAmplitudes [4362] = 8'd125;
   assign soundFileAmplitudes [4363] = 8'd124;
   assign soundFileAmplitudes [4364] = 8'd135;
   assign soundFileAmplitudes [4365] = 8'd142;
   assign soundFileAmplitudes [4366] = 8'd143;
   assign soundFileAmplitudes [4367] = 8'd152;
   assign soundFileAmplitudes [4368] = 8'd155;
   assign soundFileAmplitudes [4369] = 8'd141;
   assign soundFileAmplitudes [4370] = 8'd122;
   assign soundFileAmplitudes [4371] = 8'd109;
   assign soundFileAmplitudes [4372] = 8'd100;
   assign soundFileAmplitudes [4373] = 8'd108;
   assign soundFileAmplitudes [4374] = 8'd125;
   assign soundFileAmplitudes [4375] = 8'd137;
   assign soundFileAmplitudes [4376] = 8'd135;
   assign soundFileAmplitudes [4377] = 8'd129;
   assign soundFileAmplitudes [4378] = 8'd127;
   assign soundFileAmplitudes [4379] = 8'd135;
   assign soundFileAmplitudes [4380] = 8'd160;
   assign soundFileAmplitudes [4381] = 8'd167;
   assign soundFileAmplitudes [4382] = 8'd159;
   assign soundFileAmplitudes [4383] = 8'd142;
   assign soundFileAmplitudes [4384] = 8'd144;
   assign soundFileAmplitudes [4385] = 8'd146;
   assign soundFileAmplitudes [4386] = 8'd150;
   assign soundFileAmplitudes [4387] = 8'd162;
   assign soundFileAmplitudes [4388] = 8'd149;
   assign soundFileAmplitudes [4389] = 8'd133;
   assign soundFileAmplitudes [4390] = 8'd119;
   assign soundFileAmplitudes [4391] = 8'd110;
   assign soundFileAmplitudes [4392] = 8'd114;
   assign soundFileAmplitudes [4393] = 8'd91;
   assign soundFileAmplitudes [4394] = 8'd64;
   assign soundFileAmplitudes [4395] = 8'd75;
   assign soundFileAmplitudes [4396] = 8'd94;
   assign soundFileAmplitudes [4397] = 8'd111;
   assign soundFileAmplitudes [4398] = 8'd109;
   assign soundFileAmplitudes [4399] = 8'd97;
   assign soundFileAmplitudes [4400] = 8'd99;
   assign soundFileAmplitudes [4401] = 8'd117;
   assign soundFileAmplitudes [4402] = 8'd134;
   assign soundFileAmplitudes [4403] = 8'd147;
   assign soundFileAmplitudes [4404] = 8'd151;
   assign soundFileAmplitudes [4405] = 8'd141;
   assign soundFileAmplitudes [4406] = 8'd136;
   assign soundFileAmplitudes [4407] = 8'd133;
   assign soundFileAmplitudes [4408] = 8'd123;
   assign soundFileAmplitudes [4409] = 8'd113;
   assign soundFileAmplitudes [4410] = 8'd121;
   assign soundFileAmplitudes [4411] = 8'd122;
   assign soundFileAmplitudes [4412] = 8'd109;
   assign soundFileAmplitudes [4413] = 8'd107;
   assign soundFileAmplitudes [4414] = 8'd111;
   assign soundFileAmplitudes [4415] = 8'd119;
   assign soundFileAmplitudes [4416] = 8'd141;
   assign soundFileAmplitudes [4417] = 8'd149;
   assign soundFileAmplitudes [4418] = 8'd154;
   assign soundFileAmplitudes [4419] = 8'd159;
   assign soundFileAmplitudes [4420] = 8'd160;
   assign soundFileAmplitudes [4421] = 8'd161;
   assign soundFileAmplitudes [4422] = 8'd152;
   assign soundFileAmplitudes [4423] = 8'd139;
   assign soundFileAmplitudes [4424] = 8'd134;
   assign soundFileAmplitudes [4425] = 8'd136;
   assign soundFileAmplitudes [4426] = 8'd134;
   assign soundFileAmplitudes [4427] = 8'd123;
   assign soundFileAmplitudes [4428] = 8'd132;
   assign soundFileAmplitudes [4429] = 8'd121;
   assign soundFileAmplitudes [4430] = 8'd104;
   assign soundFileAmplitudes [4431] = 8'd102;
   assign soundFileAmplitudes [4432] = 8'd82;
   assign soundFileAmplitudes [4433] = 8'd103;
   assign soundFileAmplitudes [4434] = 8'd119;
   assign soundFileAmplitudes [4435] = 8'd116;
   assign soundFileAmplitudes [4436] = 8'd100;
   assign soundFileAmplitudes [4437] = 8'd94;
   assign soundFileAmplitudes [4438] = 8'd109;
   assign soundFileAmplitudes [4439] = 8'd128;
   assign soundFileAmplitudes [4440] = 8'd143;
   assign soundFileAmplitudes [4441] = 8'd141;
   assign soundFileAmplitudes [4442] = 8'd147;
   assign soundFileAmplitudes [4443] = 8'd140;
   assign soundFileAmplitudes [4444] = 8'd119;
   assign soundFileAmplitudes [4445] = 8'd105;
   assign soundFileAmplitudes [4446] = 8'd109;
   assign soundFileAmplitudes [4447] = 8'd111;
   assign soundFileAmplitudes [4448] = 8'd116;
   assign soundFileAmplitudes [4449] = 8'd112;
   assign soundFileAmplitudes [4450] = 8'd102;
   assign soundFileAmplitudes [4451] = 8'd101;
   assign soundFileAmplitudes [4452] = 8'd123;
   assign soundFileAmplitudes [4453] = 8'd137;
   assign soundFileAmplitudes [4454] = 8'd145;
   assign soundFileAmplitudes [4455] = 8'd142;
   assign soundFileAmplitudes [4456] = 8'd139;
   assign soundFileAmplitudes [4457] = 8'd151;
   assign soundFileAmplitudes [4458] = 8'd154;
   assign soundFileAmplitudes [4459] = 8'd158;
   assign soundFileAmplitudes [4460] = 8'd155;
   assign soundFileAmplitudes [4461] = 8'd151;
   assign soundFileAmplitudes [4462] = 8'd137;
   assign soundFileAmplitudes [4463] = 8'd137;
   assign soundFileAmplitudes [4464] = 8'd141;
   assign soundFileAmplitudes [4465] = 8'd146;
   assign soundFileAmplitudes [4466] = 8'd128;
   assign soundFileAmplitudes [4467] = 8'd125;
   assign soundFileAmplitudes [4468] = 8'd123;
   assign soundFileAmplitudes [4469] = 8'd107;
   assign soundFileAmplitudes [4470] = 8'd106;
   assign soundFileAmplitudes [4471] = 8'd82;
   assign soundFileAmplitudes [4472] = 8'd73;
   assign soundFileAmplitudes [4473] = 8'd85;
   assign soundFileAmplitudes [4474] = 8'd89;
   assign soundFileAmplitudes [4475] = 8'd95;
   assign soundFileAmplitudes [4476] = 8'd110;
   assign soundFileAmplitudes [4477] = 8'd116;
   assign soundFileAmplitudes [4478] = 8'd122;
   assign soundFileAmplitudes [4479] = 8'd120;
   assign soundFileAmplitudes [4480] = 8'd119;
   assign soundFileAmplitudes [4481] = 8'd112;
   assign soundFileAmplitudes [4482] = 8'd110;
   assign soundFileAmplitudes [4483] = 8'd114;
   assign soundFileAmplitudes [4484] = 8'd124;
   assign soundFileAmplitudes [4485] = 8'd140;
   assign soundFileAmplitudes [4486] = 8'd133;
   assign soundFileAmplitudes [4487] = 8'd130;
   assign soundFileAmplitudes [4488] = 8'd139;
   assign soundFileAmplitudes [4489] = 8'd150;
   assign soundFileAmplitudes [4490] = 8'd155;
   assign soundFileAmplitudes [4491] = 8'd153;
   assign soundFileAmplitudes [4492] = 8'd148;
   assign soundFileAmplitudes [4493] = 8'd146;
   assign soundFileAmplitudes [4494] = 8'd144;
   assign soundFileAmplitudes [4495] = 8'd149;
   assign soundFileAmplitudes [4496] = 8'd158;
   assign soundFileAmplitudes [4497] = 8'd157;
   assign soundFileAmplitudes [4498] = 8'd149;
   assign soundFileAmplitudes [4499] = 8'd140;
   assign soundFileAmplitudes [4500] = 8'd133;
   assign soundFileAmplitudes [4501] = 8'd130;
   assign soundFileAmplitudes [4502] = 8'd134;
   assign soundFileAmplitudes [4503] = 8'd131;
   assign soundFileAmplitudes [4504] = 8'd135;
   assign soundFileAmplitudes [4505] = 8'd128;
   assign soundFileAmplitudes [4506] = 8'd101;
   assign soundFileAmplitudes [4507] = 8'd115;
   assign soundFileAmplitudes [4508] = 8'd117;
   assign soundFileAmplitudes [4509] = 8'd122;
   assign soundFileAmplitudes [4510] = 8'd128;
   assign soundFileAmplitudes [4511] = 8'd87;
   assign soundFileAmplitudes [4512] = 8'd74;
   assign soundFileAmplitudes [4513] = 8'd87;
   assign soundFileAmplitudes [4514] = 8'd100;
   assign soundFileAmplitudes [4515] = 8'd100;
   assign soundFileAmplitudes [4516] = 8'd96;
   assign soundFileAmplitudes [4517] = 8'd93;
   assign soundFileAmplitudes [4518] = 8'd76;
   assign soundFileAmplitudes [4519] = 8'd80;
   assign soundFileAmplitudes [4520] = 8'd99;
   assign soundFileAmplitudes [4521] = 8'd114;
   assign soundFileAmplitudes [4522] = 8'd135;
   assign soundFileAmplitudes [4523] = 8'd152;
   assign soundFileAmplitudes [4524] = 8'd150;
   assign soundFileAmplitudes [4525] = 8'd157;
   assign soundFileAmplitudes [4526] = 8'd173;
   assign soundFileAmplitudes [4527] = 8'd154;
   assign soundFileAmplitudes [4528] = 8'd164;
   assign soundFileAmplitudes [4529] = 8'd166;
   assign soundFileAmplitudes [4530] = 8'd164;
   assign soundFileAmplitudes [4531] = 8'd179;
   assign soundFileAmplitudes [4532] = 8'd171;
   assign soundFileAmplitudes [4533] = 8'd159;
   assign soundFileAmplitudes [4534] = 8'd151;
   assign soundFileAmplitudes [4535] = 8'd153;
   assign soundFileAmplitudes [4536] = 8'd142;
   assign soundFileAmplitudes [4537] = 8'd136;
   assign soundFileAmplitudes [4538] = 8'd130;
   assign soundFileAmplitudes [4539] = 8'd131;
   assign soundFileAmplitudes [4540] = 8'd120;
   assign soundFileAmplitudes [4541] = 8'd118;
   assign soundFileAmplitudes [4542] = 8'd107;
   assign soundFileAmplitudes [4543] = 8'd94;
   assign soundFileAmplitudes [4544] = 8'd86;
   assign soundFileAmplitudes [4545] = 8'd90;
   assign soundFileAmplitudes [4546] = 8'd95;
   assign soundFileAmplitudes [4547] = 8'd100;
   assign soundFileAmplitudes [4548] = 8'd106;
   assign soundFileAmplitudes [4549] = 8'd97;
   assign soundFileAmplitudes [4550] = 8'd111;
   assign soundFileAmplitudes [4551] = 8'd103;
   assign soundFileAmplitudes [4552] = 8'd96;
   assign soundFileAmplitudes [4553] = 8'd99;
   assign soundFileAmplitudes [4554] = 8'd102;
   assign soundFileAmplitudes [4555] = 8'd88;
   assign soundFileAmplitudes [4556] = 8'd84;
   assign soundFileAmplitudes [4557] = 8'd95;
   assign soundFileAmplitudes [4558] = 8'd102;
   assign soundFileAmplitudes [4559] = 8'd123;
   assign soundFileAmplitudes [4560] = 8'd134;
   assign soundFileAmplitudes [4561] = 8'd150;
   assign soundFileAmplitudes [4562] = 8'd160;
   assign soundFileAmplitudes [4563] = 8'd171;
   assign soundFileAmplitudes [4564] = 8'd169;
   assign soundFileAmplitudes [4565] = 8'd169;
   assign soundFileAmplitudes [4566] = 8'd175;
   assign soundFileAmplitudes [4567] = 8'd173;
   assign soundFileAmplitudes [4568] = 8'd179;
   assign soundFileAmplitudes [4569] = 8'd173;
   assign soundFileAmplitudes [4570] = 8'd173;
   assign soundFileAmplitudes [4571] = 8'd162;
   assign soundFileAmplitudes [4572] = 8'd142;
   assign soundFileAmplitudes [4573] = 8'd129;
   assign soundFileAmplitudes [4574] = 8'd118;
   assign soundFileAmplitudes [4575] = 8'd108;
   assign soundFileAmplitudes [4576] = 8'd99;
   assign soundFileAmplitudes [4577] = 8'd85;
   assign soundFileAmplitudes [4578] = 8'd73;
   assign soundFileAmplitudes [4579] = 8'd73;
   assign soundFileAmplitudes [4580] = 8'd81;
   assign soundFileAmplitudes [4581] = 8'd95;
   assign soundFileAmplitudes [4582] = 8'd116;
   assign soundFileAmplitudes [4583] = 8'd134;
   assign soundFileAmplitudes [4584] = 8'd141;
   assign soundFileAmplitudes [4585] = 8'd140;
   assign soundFileAmplitudes [4586] = 8'd124;
   assign soundFileAmplitudes [4587] = 8'd114;
   assign soundFileAmplitudes [4588] = 8'd132;
   assign soundFileAmplitudes [4589] = 8'd153;
   assign soundFileAmplitudes [4590] = 8'd149;
   assign soundFileAmplitudes [4591] = 8'd130;
   assign soundFileAmplitudes [4592] = 8'd96;
   assign soundFileAmplitudes [4593] = 8'd81;
   assign soundFileAmplitudes [4594] = 8'd91;
   assign soundFileAmplitudes [4595] = 8'd87;
   assign soundFileAmplitudes [4596] = 8'd88;
   assign soundFileAmplitudes [4597] = 8'd90;
   assign soundFileAmplitudes [4598] = 8'd89;
   assign soundFileAmplitudes [4599] = 8'd100;
   assign soundFileAmplitudes [4600] = 8'd119;
   assign soundFileAmplitudes [4601] = 8'd144;
   assign soundFileAmplitudes [4602] = 8'd153;
   assign soundFileAmplitudes [4603] = 8'd163;
   assign soundFileAmplitudes [4604] = 8'd167;
   assign soundFileAmplitudes [4605] = 8'd181;
   assign soundFileAmplitudes [4606] = 8'd192;
   assign soundFileAmplitudes [4607] = 8'd187;
   assign soundFileAmplitudes [4608] = 8'd180;
   assign soundFileAmplitudes [4609] = 8'd165;
   assign soundFileAmplitudes [4610] = 8'd155;
   assign soundFileAmplitudes [4611] = 8'd145;
   assign soundFileAmplitudes [4612] = 8'd132;
   assign soundFileAmplitudes [4613] = 8'd115;
   assign soundFileAmplitudes [4614] = 8'd99;
   assign soundFileAmplitudes [4615] = 8'd86;
   assign soundFileAmplitudes [4616] = 8'd84;
   assign soundFileAmplitudes [4617] = 8'd85;
   assign soundFileAmplitudes [4618] = 8'd92;
   assign soundFileAmplitudes [4619] = 8'd97;
   assign soundFileAmplitudes [4620] = 8'd108;
   assign soundFileAmplitudes [4621] = 8'd119;
   assign soundFileAmplitudes [4622] = 8'd123;
   assign soundFileAmplitudes [4623] = 8'd122;
   assign soundFileAmplitudes [4624] = 8'd135;
   assign soundFileAmplitudes [4625] = 8'd143;
   assign soundFileAmplitudes [4626] = 8'd144;
   assign soundFileAmplitudes [4627] = 8'd136;
   assign soundFileAmplitudes [4628] = 8'd116;
   assign soundFileAmplitudes [4629] = 8'd94;
   assign soundFileAmplitudes [4630] = 8'd88;
   assign soundFileAmplitudes [4631] = 8'd91;
   assign soundFileAmplitudes [4632] = 8'd96;
   assign soundFileAmplitudes [4633] = 8'd107;
   assign soundFileAmplitudes [4634] = 8'd105;
   assign soundFileAmplitudes [4635] = 8'd108;
   assign soundFileAmplitudes [4636] = 8'd112;
   assign soundFileAmplitudes [4637] = 8'd119;
   assign soundFileAmplitudes [4638] = 8'd126;
   assign soundFileAmplitudes [4639] = 8'd137;
   assign soundFileAmplitudes [4640] = 8'd140;
   assign soundFileAmplitudes [4641] = 8'd155;
   assign soundFileAmplitudes [4642] = 8'd160;
   assign soundFileAmplitudes [4643] = 8'd170;
   assign soundFileAmplitudes [4644] = 8'd184;
   assign soundFileAmplitudes [4645] = 8'd167;
   assign soundFileAmplitudes [4646] = 8'd168;
   assign soundFileAmplitudes [4647] = 8'd163;
   assign soundFileAmplitudes [4648] = 8'd165;
   assign soundFileAmplitudes [4649] = 8'd154;
   assign soundFileAmplitudes [4650] = 8'd133;
   assign soundFileAmplitudes [4651] = 8'd122;
   assign soundFileAmplitudes [4652] = 8'd101;
   assign soundFileAmplitudes [4653] = 8'd86;
   assign soundFileAmplitudes [4654] = 8'd81;
   assign soundFileAmplitudes [4655] = 8'd86;
   assign soundFileAmplitudes [4656] = 8'd103;
   assign soundFileAmplitudes [4657] = 8'd125;
   assign soundFileAmplitudes [4658] = 8'd122;
   assign soundFileAmplitudes [4659] = 8'd113;
   assign soundFileAmplitudes [4660] = 8'd115;
   assign soundFileAmplitudes [4661] = 8'd132;
   assign soundFileAmplitudes [4662] = 8'd151;
   assign soundFileAmplitudes [4663] = 8'd153;
   assign soundFileAmplitudes [4664] = 8'd165;
   assign soundFileAmplitudes [4665] = 8'd154;
   assign soundFileAmplitudes [4666] = 8'd134;
   assign soundFileAmplitudes [4667] = 8'd111;
   assign soundFileAmplitudes [4668] = 8'd98;
   assign soundFileAmplitudes [4669] = 8'd102;
   assign soundFileAmplitudes [4670] = 8'd104;
   assign soundFileAmplitudes [4671] = 8'd101;
   assign soundFileAmplitudes [4672] = 8'd90;
   assign soundFileAmplitudes [4673] = 8'd98;
   assign soundFileAmplitudes [4674] = 8'd112;
   assign soundFileAmplitudes [4675] = 8'd109;
   assign soundFileAmplitudes [4676] = 8'd124;
   assign soundFileAmplitudes [4677] = 8'd137;
   assign soundFileAmplitudes [4678] = 8'd129;
   assign soundFileAmplitudes [4679] = 8'd144;
   assign soundFileAmplitudes [4680] = 8'd138;
   assign soundFileAmplitudes [4681] = 8'd155;
   assign soundFileAmplitudes [4682] = 8'd165;
   assign soundFileAmplitudes [4683] = 8'd144;
   assign soundFileAmplitudes [4684] = 8'd132;
   assign soundFileAmplitudes [4685] = 8'd125;
   assign soundFileAmplitudes [4686] = 8'd133;
   assign soundFileAmplitudes [4687] = 8'd134;
   assign soundFileAmplitudes [4688] = 8'd131;
   assign soundFileAmplitudes [4689] = 8'd125;
   assign soundFileAmplitudes [4690] = 8'd109;
   assign soundFileAmplitudes [4691] = 8'd103;
   assign soundFileAmplitudes [4692] = 8'd110;
   assign soundFileAmplitudes [4693] = 8'd104;
   assign soundFileAmplitudes [4694] = 8'd110;
   assign soundFileAmplitudes [4695] = 8'd114;
   assign soundFileAmplitudes [4696] = 8'd106;
   assign soundFileAmplitudes [4697] = 8'd123;
   assign soundFileAmplitudes [4698] = 8'd146;
   assign soundFileAmplitudes [4699] = 8'd156;
   assign soundFileAmplitudes [4700] = 8'd174;
   assign soundFileAmplitudes [4701] = 8'd168;
   assign soundFileAmplitudes [4702] = 8'd138;
   assign soundFileAmplitudes [4703] = 8'd114;
   assign soundFileAmplitudes [4704] = 8'd91;
   assign soundFileAmplitudes [4705] = 8'd84;
   assign soundFileAmplitudes [4706] = 8'd104;
   assign soundFileAmplitudes [4707] = 8'd122;
   assign soundFileAmplitudes [4708] = 8'd112;
   assign soundFileAmplitudes [4709] = 8'd111;
   assign soundFileAmplitudes [4710] = 8'd106;
   assign soundFileAmplitudes [4711] = 8'd94;
   assign soundFileAmplitudes [4712] = 8'd105;
   assign soundFileAmplitudes [4713] = 8'd120;
   assign soundFileAmplitudes [4714] = 8'd139;
   assign soundFileAmplitudes [4715] = 8'd148;
   assign soundFileAmplitudes [4716] = 8'd147;
   assign soundFileAmplitudes [4717] = 8'd146;
   assign soundFileAmplitudes [4718] = 8'd127;
   assign soundFileAmplitudes [4719] = 8'd125;
   assign soundFileAmplitudes [4720] = 8'd118;
   assign soundFileAmplitudes [4721] = 8'd116;
   assign soundFileAmplitudes [4722] = 8'd128;
   assign soundFileAmplitudes [4723] = 8'd143;
   assign soundFileAmplitudes [4724] = 8'd154;
   assign soundFileAmplitudes [4725] = 8'd135;
   assign soundFileAmplitudes [4726] = 8'd125;
   assign soundFileAmplitudes [4727] = 8'd113;
   assign soundFileAmplitudes [4728] = 8'd108;
   assign soundFileAmplitudes [4729] = 8'd119;
   assign soundFileAmplitudes [4730] = 8'd133;
   assign soundFileAmplitudes [4731] = 8'd148;
   assign soundFileAmplitudes [4732] = 8'd141;
   assign soundFileAmplitudes [4733] = 8'd127;
   assign soundFileAmplitudes [4734] = 8'd133;
   assign soundFileAmplitudes [4735] = 8'd146;
   assign soundFileAmplitudes [4736] = 8'd138;
   assign soundFileAmplitudes [4737] = 8'd142;
   assign soundFileAmplitudes [4738] = 8'd136;
   assign soundFileAmplitudes [4739] = 8'd129;
   assign soundFileAmplitudes [4740] = 8'd112;
   assign soundFileAmplitudes [4741] = 8'd98;
   assign soundFileAmplitudes [4742] = 8'd114;
   assign soundFileAmplitudes [4743] = 8'd112;
   assign soundFileAmplitudes [4744] = 8'd119;
   assign soundFileAmplitudes [4745] = 8'd113;
   assign soundFileAmplitudes [4746] = 8'd116;
   assign soundFileAmplitudes [4747] = 8'd119;
   assign soundFileAmplitudes [4748] = 8'd118;
   assign soundFileAmplitudes [4749] = 8'd124;
   assign soundFileAmplitudes [4750] = 8'd122;
   assign soundFileAmplitudes [4751] = 8'd120;
   assign soundFileAmplitudes [4752] = 8'd132;
   assign soundFileAmplitudes [4753] = 8'd136;
   assign soundFileAmplitudes [4754] = 8'd120;
   assign soundFileAmplitudes [4755] = 8'd128;
   assign soundFileAmplitudes [4756] = 8'd117;
   assign soundFileAmplitudes [4757] = 8'd116;
   assign soundFileAmplitudes [4758] = 8'd112;
   assign soundFileAmplitudes [4759] = 8'd106;
   assign soundFileAmplitudes [4760] = 8'd111;
   assign soundFileAmplitudes [4761] = 8'd106;
   assign soundFileAmplitudes [4762] = 8'd117;
   assign soundFileAmplitudes [4763] = 8'd112;
   assign soundFileAmplitudes [4764] = 8'd118;
   assign soundFileAmplitudes [4765] = 8'd121;
   assign soundFileAmplitudes [4766] = 8'd121;
   assign soundFileAmplitudes [4767] = 8'd132;
   assign soundFileAmplitudes [4768] = 8'd136;
   assign soundFileAmplitudes [4769] = 8'd137;
   assign soundFileAmplitudes [4770] = 8'd166;
   assign soundFileAmplitudes [4771] = 8'd177;
   assign soundFileAmplitudes [4772] = 8'd167;
   assign soundFileAmplitudes [4773] = 8'd168;
   assign soundFileAmplitudes [4774] = 8'd146;
   assign soundFileAmplitudes [4775] = 8'd132;
   assign soundFileAmplitudes [4776] = 8'd130;
   assign soundFileAmplitudes [4777] = 8'd134;
   assign soundFileAmplitudes [4778] = 8'd131;
   assign soundFileAmplitudes [4779] = 8'd130;
   assign soundFileAmplitudes [4780] = 8'd121;
   assign soundFileAmplitudes [4781] = 8'd109;
   assign soundFileAmplitudes [4782] = 8'd112;
   assign soundFileAmplitudes [4783] = 8'd107;
   assign soundFileAmplitudes [4784] = 8'd113;
   assign soundFileAmplitudes [4785] = 8'd117;
   assign soundFileAmplitudes [4786] = 8'd126;
   assign soundFileAmplitudes [4787] = 8'd134;
   assign soundFileAmplitudes [4788] = 8'd132;
   assign soundFileAmplitudes [4789] = 8'd109;
   assign soundFileAmplitudes [4790] = 8'd105;
   assign soundFileAmplitudes [4791] = 8'd104;
   assign soundFileAmplitudes [4792] = 8'd105;
   assign soundFileAmplitudes [4793] = 8'd123;
   assign soundFileAmplitudes [4794] = 8'd123;
   assign soundFileAmplitudes [4795] = 8'd125;
   assign soundFileAmplitudes [4796] = 8'd110;
   assign soundFileAmplitudes [4797] = 8'd99;
   assign soundFileAmplitudes [4798] = 8'd94;
   assign soundFileAmplitudes [4799] = 8'd95;
   assign soundFileAmplitudes [4800] = 8'd119;
   assign soundFileAmplitudes [4801] = 8'd137;
   assign soundFileAmplitudes [4802] = 8'd146;
   assign soundFileAmplitudes [4803] = 8'd149;
   assign soundFileAmplitudes [4804] = 8'd143;
   assign soundFileAmplitudes [4805] = 8'd141;
   assign soundFileAmplitudes [4806] = 8'd153;
   assign soundFileAmplitudes [4807] = 8'd171;
   assign soundFileAmplitudes [4808] = 8'd169;
   assign soundFileAmplitudes [4809] = 8'd165;
   assign soundFileAmplitudes [4810] = 8'd151;
   assign soundFileAmplitudes [4811] = 8'd139;
   assign soundFileAmplitudes [4812] = 8'd138;
   assign soundFileAmplitudes [4813] = 8'd129;
   assign soundFileAmplitudes [4814] = 8'd121;
   assign soundFileAmplitudes [4815] = 8'd110;
   assign soundFileAmplitudes [4816] = 8'd97;
   assign soundFileAmplitudes [4817] = 8'd96;
   assign soundFileAmplitudes [4818] = 8'd86;
   assign soundFileAmplitudes [4819] = 8'd88;
   assign soundFileAmplitudes [4820] = 8'd109;
   assign soundFileAmplitudes [4821] = 8'd120;
   assign soundFileAmplitudes [4822] = 8'd142;
   assign soundFileAmplitudes [4823] = 8'd146;
   assign soundFileAmplitudes [4824] = 8'd137;
   assign soundFileAmplitudes [4825] = 8'd123;
   assign soundFileAmplitudes [4826] = 8'd124;
   assign soundFileAmplitudes [4827] = 8'd129;
   assign soundFileAmplitudes [4828] = 8'd139;
   assign soundFileAmplitudes [4829] = 8'd129;
   assign soundFileAmplitudes [4830] = 8'd111;
   assign soundFileAmplitudes [4831] = 8'd97;
   assign soundFileAmplitudes [4832] = 8'd110;
   assign soundFileAmplitudes [4833] = 8'd127;
   assign soundFileAmplitudes [4834] = 8'd101;
   assign soundFileAmplitudes [4835] = 8'd103;
   assign soundFileAmplitudes [4836] = 8'd115;
   assign soundFileAmplitudes [4837] = 8'd138;
   assign soundFileAmplitudes [4838] = 8'd142;
   assign soundFileAmplitudes [4839] = 8'd139;
   assign soundFileAmplitudes [4840] = 8'd138;
   assign soundFileAmplitudes [4841] = 8'd137;
   assign soundFileAmplitudes [4842] = 8'd151;
   assign soundFileAmplitudes [4843] = 8'd160;
   assign soundFileAmplitudes [4844] = 8'd156;
   assign soundFileAmplitudes [4845] = 8'd147;
   assign soundFileAmplitudes [4846] = 8'd129;
   assign soundFileAmplitudes [4847] = 8'd114;
   assign soundFileAmplitudes [4848] = 8'd121;
   assign soundFileAmplitudes [4849] = 8'd122;
   assign soundFileAmplitudes [4850] = 8'd119;
   assign soundFileAmplitudes [4851] = 8'd122;
   assign soundFileAmplitudes [4852] = 8'd114;
   assign soundFileAmplitudes [4853] = 8'd96;
   assign soundFileAmplitudes [4854] = 8'd83;
   assign soundFileAmplitudes [4855] = 8'd79;
   assign soundFileAmplitudes [4856] = 8'd75;
   assign soundFileAmplitudes [4857] = 8'd85;
   assign soundFileAmplitudes [4858] = 8'd110;
   assign soundFileAmplitudes [4859] = 8'd119;
   assign soundFileAmplitudes [4860] = 8'd126;
   assign soundFileAmplitudes [4861] = 8'd138;
   assign soundFileAmplitudes [4862] = 8'd136;
   assign soundFileAmplitudes [4863] = 8'd127;
   assign soundFileAmplitudes [4864] = 8'd133;
   assign soundFileAmplitudes [4865] = 8'd148;
   assign soundFileAmplitudes [4866] = 8'd148;
   assign soundFileAmplitudes [4867] = 8'd135;
   assign soundFileAmplitudes [4868] = 8'd141;
   assign soundFileAmplitudes [4869] = 8'd139;
   assign soundFileAmplitudes [4870] = 8'd140;
   assign soundFileAmplitudes [4871] = 8'd131;
   assign soundFileAmplitudes [4872] = 8'd130;
   assign soundFileAmplitudes [4873] = 8'd152;
   assign soundFileAmplitudes [4874] = 8'd161;
   assign soundFileAmplitudes [4875] = 8'd168;
   assign soundFileAmplitudes [4876] = 8'd161;
   assign soundFileAmplitudes [4877] = 8'd146;
   assign soundFileAmplitudes [4878] = 8'd127;
   assign soundFileAmplitudes [4879] = 8'd129;
   assign soundFileAmplitudes [4880] = 8'd125;
   assign soundFileAmplitudes [4881] = 8'd120;
   assign soundFileAmplitudes [4882] = 8'd127;
   assign soundFileAmplitudes [4883] = 8'd137;
   assign soundFileAmplitudes [4884] = 8'd143;
   assign soundFileAmplitudes [4885] = 8'd125;
   assign soundFileAmplitudes [4886] = 8'd120;
   assign soundFileAmplitudes [4887] = 8'd107;
   assign soundFileAmplitudes [4888] = 8'd101;
   assign soundFileAmplitudes [4889] = 8'd97;
   assign soundFileAmplitudes [4890] = 8'd84;
   assign soundFileAmplitudes [4891] = 8'd81;
   assign soundFileAmplitudes [4892] = 8'd73;
   assign soundFileAmplitudes [4893] = 8'd77;
   assign soundFileAmplitudes [4894] = 8'd81;
   assign soundFileAmplitudes [4895] = 8'd78;
   assign soundFileAmplitudes [4896] = 8'd85;
   assign soundFileAmplitudes [4897] = 8'd96;
   assign soundFileAmplitudes [4898] = 8'd111;
   assign soundFileAmplitudes [4899] = 8'd128;
   assign soundFileAmplitudes [4900] = 8'd144;
   assign soundFileAmplitudes [4901] = 8'd152;
   assign soundFileAmplitudes [4902] = 8'd152;
   assign soundFileAmplitudes [4903] = 8'd160;
   assign soundFileAmplitudes [4904] = 8'd160;
   assign soundFileAmplitudes [4905] = 8'd163;
   assign soundFileAmplitudes [4906] = 8'd160;
   assign soundFileAmplitudes [4907] = 8'd162;
   assign soundFileAmplitudes [4908] = 8'd162;
   assign soundFileAmplitudes [4909] = 8'd152;
   assign soundFileAmplitudes [4910] = 8'd151;
   assign soundFileAmplitudes [4911] = 8'd163;
   assign soundFileAmplitudes [4912] = 8'd169;
   assign soundFileAmplitudes [4913] = 8'd146;
   assign soundFileAmplitudes [4914] = 8'd142;
   assign soundFileAmplitudes [4915] = 8'd150;
   assign soundFileAmplitudes [4916] = 8'd141;
   assign soundFileAmplitudes [4917] = 8'd120;
   assign soundFileAmplitudes [4918] = 8'd118;
   assign soundFileAmplitudes [4919] = 8'd118;
   assign soundFileAmplitudes [4920] = 8'd118;
   assign soundFileAmplitudes [4921] = 8'd111;
   assign soundFileAmplitudes [4922] = 8'd96;
   assign soundFileAmplitudes [4923] = 8'd93;
   assign soundFileAmplitudes [4924] = 8'd93;
   assign soundFileAmplitudes [4925] = 8'd101;
   assign soundFileAmplitudes [4926] = 8'd110;
   assign soundFileAmplitudes [4927] = 8'd105;
   assign soundFileAmplitudes [4928] = 8'd94;
   assign soundFileAmplitudes [4929] = 8'd87;
   assign soundFileAmplitudes [4930] = 8'd83;
   assign soundFileAmplitudes [4931] = 8'd85;
   assign soundFileAmplitudes [4932] = 8'd97;
   assign soundFileAmplitudes [4933] = 8'd111;
   assign soundFileAmplitudes [4934] = 8'd114;
   assign soundFileAmplitudes [4935] = 8'd125;
   assign soundFileAmplitudes [4936] = 8'd125;
   assign soundFileAmplitudes [4937] = 8'd122;
   assign soundFileAmplitudes [4938] = 8'd133;
   assign soundFileAmplitudes [4939] = 8'd120;
   assign soundFileAmplitudes [4940] = 8'd130;
   assign soundFileAmplitudes [4941] = 8'd145;
   assign soundFileAmplitudes [4942] = 8'd142;
   assign soundFileAmplitudes [4943] = 8'd143;
   assign soundFileAmplitudes [4944] = 8'd143;
   assign soundFileAmplitudes [4945] = 8'd152;
   assign soundFileAmplitudes [4946] = 8'd159;
   assign soundFileAmplitudes [4947] = 8'd169;
   assign soundFileAmplitudes [4948] = 8'd162;
   assign soundFileAmplitudes [4949] = 8'd170;
   assign soundFileAmplitudes [4950] = 8'd170;
   assign soundFileAmplitudes [4951] = 8'd166;
   assign soundFileAmplitudes [4952] = 8'd160;
   assign soundFileAmplitudes [4953] = 8'd149;
   assign soundFileAmplitudes [4954] = 8'd147;
   assign soundFileAmplitudes [4955] = 8'd123;
   assign soundFileAmplitudes [4956] = 8'd121;
   assign soundFileAmplitudes [4957] = 8'd110;
   assign soundFileAmplitudes [4958] = 8'd110;
   assign soundFileAmplitudes [4959] = 8'd117;
   assign soundFileAmplitudes [4960] = 8'd118;
   assign soundFileAmplitudes [4961] = 8'd120;
   assign soundFileAmplitudes [4962] = 8'd116;
   assign soundFileAmplitudes [4963] = 8'd120;
   assign soundFileAmplitudes [4964] = 8'd113;
   assign soundFileAmplitudes [4965] = 8'd101;
   assign soundFileAmplitudes [4966] = 8'd86;
   assign soundFileAmplitudes [4967] = 8'd79;
   assign soundFileAmplitudes [4968] = 8'd84;
   assign soundFileAmplitudes [4969] = 8'd95;
   assign soundFileAmplitudes [4970] = 8'd100;
   assign soundFileAmplitudes [4971] = 8'd103;
   assign soundFileAmplitudes [4972] = 8'd113;
   assign soundFileAmplitudes [4973] = 8'd123;
   assign soundFileAmplitudes [4974] = 8'd121;
   assign soundFileAmplitudes [4975] = 8'd116;
   assign soundFileAmplitudes [4976] = 8'd115;
   assign soundFileAmplitudes [4977] = 8'd123;
   assign soundFileAmplitudes [4978] = 8'd129;
   assign soundFileAmplitudes [4979] = 8'd119;
   assign soundFileAmplitudes [4980] = 8'd118;
   assign soundFileAmplitudes [4981] = 8'd128;
   assign soundFileAmplitudes [4982] = 8'd139;
   assign soundFileAmplitudes [4983] = 8'd139;
   assign soundFileAmplitudes [4984] = 8'd137;
   assign soundFileAmplitudes [4985] = 8'd135;
   assign soundFileAmplitudes [4986] = 8'd140;
   assign soundFileAmplitudes [4987] = 8'd147;
   assign soundFileAmplitudes [4988] = 8'd162;
   assign soundFileAmplitudes [4989] = 8'd175;
   assign soundFileAmplitudes [4990] = 8'd166;
   assign soundFileAmplitudes [4991] = 8'd162;
   assign soundFileAmplitudes [4992] = 8'd150;
   assign soundFileAmplitudes [4993] = 8'd133;
   assign soundFileAmplitudes [4994] = 8'd127;
   assign soundFileAmplitudes [4995] = 8'd125;
   assign soundFileAmplitudes [4996] = 8'd129;
   assign soundFileAmplitudes [4997] = 8'd133;
   assign soundFileAmplitudes [4998] = 8'd129;
   assign soundFileAmplitudes [4999] = 8'd122;
   assign soundFileAmplitudes [5000] = 8'd114;
   assign soundFileAmplitudes [5001] = 8'd112;
   assign soundFileAmplitudes [5002] = 8'd104;
   assign soundFileAmplitudes [5003] = 8'd103;
   assign soundFileAmplitudes [5004] = 8'd101;
   assign soundFileAmplitudes [5005] = 8'd97;
   assign soundFileAmplitudes [5006] = 8'd100;
   assign soundFileAmplitudes [5007] = 8'd92;
   assign soundFileAmplitudes [5008] = 8'd83;
   assign soundFileAmplitudes [5009] = 8'd84;
   assign soundFileAmplitudes [5010] = 8'd102;
   assign soundFileAmplitudes [5011] = 8'd117;
   assign soundFileAmplitudes [5012] = 8'd123;
   assign soundFileAmplitudes [5013] = 8'd121;
   assign soundFileAmplitudes [5014] = 8'd114;
   assign soundFileAmplitudes [5015] = 8'd117;
   assign soundFileAmplitudes [5016] = 8'd117;
   assign soundFileAmplitudes [5017] = 8'd133;
   assign soundFileAmplitudes [5018] = 8'd147;
   assign soundFileAmplitudes [5019] = 8'd154;
   assign soundFileAmplitudes [5020] = 8'd156;
   assign soundFileAmplitudes [5021] = 8'd148;
   assign soundFileAmplitudes [5022] = 8'd133;
   assign soundFileAmplitudes [5023] = 8'd131;
   assign soundFileAmplitudes [5024] = 8'd143;
   assign soundFileAmplitudes [5025] = 8'd149;
   assign soundFileAmplitudes [5026] = 8'd145;
   assign soundFileAmplitudes [5027] = 8'd136;
   assign soundFileAmplitudes [5028] = 8'd125;
   assign soundFileAmplitudes [5029] = 8'd132;
   assign soundFileAmplitudes [5030] = 8'd138;
   assign soundFileAmplitudes [5031] = 8'd129;
   assign soundFileAmplitudes [5032] = 8'd144;
   assign soundFileAmplitudes [5033] = 8'd144;
   assign soundFileAmplitudes [5034] = 8'd143;
   assign soundFileAmplitudes [5035] = 8'd137;
   assign soundFileAmplitudes [5036] = 8'd130;
   assign soundFileAmplitudes [5037] = 8'd127;
   assign soundFileAmplitudes [5038] = 8'd124;
   assign soundFileAmplitudes [5039] = 8'd133;
   assign soundFileAmplitudes [5040] = 8'd127;
   assign soundFileAmplitudes [5041] = 8'd119;
   assign soundFileAmplitudes [5042] = 8'd100;
   assign soundFileAmplitudes [5043] = 8'd86;
   assign soundFileAmplitudes [5044] = 8'd86;
   assign soundFileAmplitudes [5045] = 8'd98;
   assign soundFileAmplitudes [5046] = 8'd112;
   assign soundFileAmplitudes [5047] = 8'd126;
   assign soundFileAmplitudes [5048] = 8'd127;
   assign soundFileAmplitudes [5049] = 8'd120;
   assign soundFileAmplitudes [5050] = 8'd114;
   assign soundFileAmplitudes [5051] = 8'd113;
   assign soundFileAmplitudes [5052] = 8'd116;
   assign soundFileAmplitudes [5053] = 8'd118;
   assign soundFileAmplitudes [5054] = 8'd130;
   assign soundFileAmplitudes [5055] = 8'd131;
   assign soundFileAmplitudes [5056] = 8'd128;
   assign soundFileAmplitudes [5057] = 8'd124;
   assign soundFileAmplitudes [5058] = 8'd119;
   assign soundFileAmplitudes [5059] = 8'd125;
   assign soundFileAmplitudes [5060] = 8'd137;
   assign soundFileAmplitudes [5061] = 8'd146;
   assign soundFileAmplitudes [5062] = 8'd152;
   assign soundFileAmplitudes [5063] = 8'd149;
   assign soundFileAmplitudes [5064] = 8'd154;
   assign soundFileAmplitudes [5065] = 8'd148;
   assign soundFileAmplitudes [5066] = 8'd147;
   assign soundFileAmplitudes [5067] = 8'd149;
   assign soundFileAmplitudes [5068] = 8'd134;
   assign soundFileAmplitudes [5069] = 8'd130;
   assign soundFileAmplitudes [5070] = 8'd125;
   assign soundFileAmplitudes [5071] = 8'd124;
   assign soundFileAmplitudes [5072] = 8'd124;
   assign soundFileAmplitudes [5073] = 8'd117;
   assign soundFileAmplitudes [5074] = 8'd111;
   assign soundFileAmplitudes [5075] = 8'd121;
   assign soundFileAmplitudes [5076] = 8'd124;
   assign soundFileAmplitudes [5077] = 8'd116;
   assign soundFileAmplitudes [5078] = 8'd114;
   assign soundFileAmplitudes [5079] = 8'd95;
   assign soundFileAmplitudes [5080] = 8'd89;
   assign soundFileAmplitudes [5081] = 8'd96;
   assign soundFileAmplitudes [5082] = 8'd108;
   assign soundFileAmplitudes [5083] = 8'd117;
   assign soundFileAmplitudes [5084] = 8'd118;
   assign soundFileAmplitudes [5085] = 8'd127;
   assign soundFileAmplitudes [5086] = 8'd129;
   assign soundFileAmplitudes [5087] = 8'd140;
   assign soundFileAmplitudes [5088] = 8'd145;
   assign soundFileAmplitudes [5089] = 8'd137;
   assign soundFileAmplitudes [5090] = 8'd137;
   assign soundFileAmplitudes [5091] = 8'd142;
   assign soundFileAmplitudes [5092] = 8'd142;
   assign soundFileAmplitudes [5093] = 8'd142;
   assign soundFileAmplitudes [5094] = 8'd145;
   assign soundFileAmplitudes [5095] = 8'd135;
   assign soundFileAmplitudes [5096] = 8'd124;
   assign soundFileAmplitudes [5097] = 8'd121;
   assign soundFileAmplitudes [5098] = 8'd127;
   assign soundFileAmplitudes [5099] = 8'd123;
   assign soundFileAmplitudes [5100] = 8'd119;
   assign soundFileAmplitudes [5101] = 8'd117;
   assign soundFileAmplitudes [5102] = 8'd125;
   assign soundFileAmplitudes [5103] = 8'd138;
   assign soundFileAmplitudes [5104] = 8'd131;
   assign soundFileAmplitudes [5105] = 8'd128;
   assign soundFileAmplitudes [5106] = 8'd127;
   assign soundFileAmplitudes [5107] = 8'd123;
   assign soundFileAmplitudes [5108] = 8'd125;
   assign soundFileAmplitudes [5109] = 8'd131;
   assign soundFileAmplitudes [5110] = 8'd124;
   assign soundFileAmplitudes [5111] = 8'd115;
   assign soundFileAmplitudes [5112] = 8'd110;
   assign soundFileAmplitudes [5113] = 8'd106;
   assign soundFileAmplitudes [5114] = 8'd106;
   assign soundFileAmplitudes [5115] = 8'd105;
   assign soundFileAmplitudes [5116] = 8'd114;
   assign soundFileAmplitudes [5117] = 8'd120;
   assign soundFileAmplitudes [5118] = 8'd120;
   assign soundFileAmplitudes [5119] = 8'd122;
   assign soundFileAmplitudes [5120] = 8'd134;
   assign soundFileAmplitudes [5121] = 8'd136;
   assign soundFileAmplitudes [5122] = 8'd137;
   assign soundFileAmplitudes [5123] = 8'd137;
   assign soundFileAmplitudes [5124] = 8'd129;
   assign soundFileAmplitudes [5125] = 8'd125;
   assign soundFileAmplitudes [5126] = 8'd113;
   assign soundFileAmplitudes [5127] = 8'd120;
   assign soundFileAmplitudes [5128] = 8'd132;
   assign soundFileAmplitudes [5129] = 8'd141;
   assign soundFileAmplitudes [5130] = 8'd150;
   assign soundFileAmplitudes [5131] = 8'd135;
   assign soundFileAmplitudes [5132] = 8'd124;
   assign soundFileAmplitudes [5133] = 8'd119;
   assign soundFileAmplitudes [5134] = 8'd129;
   assign soundFileAmplitudes [5135] = 8'd150;
   assign soundFileAmplitudes [5136] = 8'd149;
   assign soundFileAmplitudes [5137] = 8'd143;
   assign soundFileAmplitudes [5138] = 8'd133;
   assign soundFileAmplitudes [5139] = 8'd114;
   assign soundFileAmplitudes [5140] = 8'd108;
   assign soundFileAmplitudes [5141] = 8'd108;
   assign soundFileAmplitudes [5142] = 8'd100;
   assign soundFileAmplitudes [5143] = 8'd102;
   assign soundFileAmplitudes [5144] = 8'd106;
   assign soundFileAmplitudes [5145] = 8'd112;
   assign soundFileAmplitudes [5146] = 8'd119;
   assign soundFileAmplitudes [5147] = 8'd111;
   assign soundFileAmplitudes [5148] = 8'd105;
   assign soundFileAmplitudes [5149] = 8'd102;
   assign soundFileAmplitudes [5150] = 8'd116;
   assign soundFileAmplitudes [5151] = 8'd132;
   assign soundFileAmplitudes [5152] = 8'd136;
   assign soundFileAmplitudes [5153] = 8'd135;
   assign soundFileAmplitudes [5154] = 8'd129;
   assign soundFileAmplitudes [5155] = 8'd130;
   assign soundFileAmplitudes [5156] = 8'd128;
   assign soundFileAmplitudes [5157] = 8'd130;
   assign soundFileAmplitudes [5158] = 8'd137;
   assign soundFileAmplitudes [5159] = 8'd131;
   assign soundFileAmplitudes [5160] = 8'd127;
   assign soundFileAmplitudes [5161] = 8'd124;
   assign soundFileAmplitudes [5162] = 8'd130;
   assign soundFileAmplitudes [5163] = 8'd132;
   assign soundFileAmplitudes [5164] = 8'd142;
   assign soundFileAmplitudes [5165] = 8'd145;
   assign soundFileAmplitudes [5166] = 8'd150;
   assign soundFileAmplitudes [5167] = 8'd149;
   assign soundFileAmplitudes [5168] = 8'd128;
   assign soundFileAmplitudes [5169] = 8'd124;
   assign soundFileAmplitudes [5170] = 8'd122;
   assign soundFileAmplitudes [5171] = 8'd128;
   assign soundFileAmplitudes [5172] = 8'd137;
   assign soundFileAmplitudes [5173] = 8'd139;
   assign soundFileAmplitudes [5174] = 8'd124;
   assign soundFileAmplitudes [5175] = 8'd120;
   assign soundFileAmplitudes [5176] = 8'd126;
   assign soundFileAmplitudes [5177] = 8'd133;
   assign soundFileAmplitudes [5178] = 8'd125;
   assign soundFileAmplitudes [5179] = 8'd109;
   assign soundFileAmplitudes [5180] = 8'd106;
   assign soundFileAmplitudes [5181] = 8'd101;
   assign soundFileAmplitudes [5182] = 8'd108;
   assign soundFileAmplitudes [5183] = 8'd111;
   assign soundFileAmplitudes [5184] = 8'd102;
   assign soundFileAmplitudes [5185] = 8'd104;
   assign soundFileAmplitudes [5186] = 8'd108;
   assign soundFileAmplitudes [5187] = 8'd111;
   assign soundFileAmplitudes [5188] = 8'd116;
   assign soundFileAmplitudes [5189] = 8'd120;
   assign soundFileAmplitudes [5190] = 8'd138;
   assign soundFileAmplitudes [5191] = 8'd148;
   assign soundFileAmplitudes [5192] = 8'd154;
   assign soundFileAmplitudes [5193] = 8'd153;
   assign soundFileAmplitudes [5194] = 8'd142;
   assign soundFileAmplitudes [5195] = 8'd137;
   assign soundFileAmplitudes [5196] = 8'd142;
   assign soundFileAmplitudes [5197] = 8'd154;
   assign soundFileAmplitudes [5198] = 8'd160;
   assign soundFileAmplitudes [5199] = 8'd148;
   assign soundFileAmplitudes [5200] = 8'd134;
   assign soundFileAmplitudes [5201] = 8'd120;
   assign soundFileAmplitudes [5202] = 8'd116;
   assign soundFileAmplitudes [5203] = 8'd130;
   assign soundFileAmplitudes [5204] = 8'd123;
   assign soundFileAmplitudes [5205] = 8'd111;
   assign soundFileAmplitudes [5206] = 8'd112;
   assign soundFileAmplitudes [5207] = 8'd112;
   assign soundFileAmplitudes [5208] = 8'd107;
   assign soundFileAmplitudes [5209] = 8'd103;
   assign soundFileAmplitudes [5210] = 8'd110;
   assign soundFileAmplitudes [5211] = 8'd122;
   assign soundFileAmplitudes [5212] = 8'd127;
   assign soundFileAmplitudes [5213] = 8'd135;
   assign soundFileAmplitudes [5214] = 8'd137;
   assign soundFileAmplitudes [5215] = 8'd138;
   assign soundFileAmplitudes [5216] = 8'd114;
   assign soundFileAmplitudes [5217] = 8'd104;
   assign soundFileAmplitudes [5218] = 8'd114;
   assign soundFileAmplitudes [5219] = 8'd125;
   assign soundFileAmplitudes [5220] = 8'd141;
   assign soundFileAmplitudes [5221] = 8'd138;
   assign soundFileAmplitudes [5222] = 8'd124;
   assign soundFileAmplitudes [5223] = 8'd107;
   assign soundFileAmplitudes [5224] = 8'd104;
   assign soundFileAmplitudes [5225] = 8'd116;
   assign soundFileAmplitudes [5226] = 8'd135;
   assign soundFileAmplitudes [5227] = 8'd142;
   assign soundFileAmplitudes [5228] = 8'd147;
   assign soundFileAmplitudes [5229] = 8'd147;
   assign soundFileAmplitudes [5230] = 8'd144;
   assign soundFileAmplitudes [5231] = 8'd141;
   assign soundFileAmplitudes [5232] = 8'd149;
   assign soundFileAmplitudes [5233] = 8'd154;
   assign soundFileAmplitudes [5234] = 8'd153;
   assign soundFileAmplitudes [5235] = 8'd143;
   assign soundFileAmplitudes [5236] = 8'd125;
   assign soundFileAmplitudes [5237] = 8'd116;
   assign soundFileAmplitudes [5238] = 8'd101;
   assign soundFileAmplitudes [5239] = 8'd106;
   assign soundFileAmplitudes [5240] = 8'd101;
   assign soundFileAmplitudes [5241] = 8'd100;
   assign soundFileAmplitudes [5242] = 8'd104;
   assign soundFileAmplitudes [5243] = 8'd113;
   assign soundFileAmplitudes [5244] = 8'd113;
   assign soundFileAmplitudes [5245] = 8'd109;
   assign soundFileAmplitudes [5246] = 8'd108;
   assign soundFileAmplitudes [5247] = 8'd109;
   assign soundFileAmplitudes [5248] = 8'd128;
   assign soundFileAmplitudes [5249] = 8'd143;
   assign soundFileAmplitudes [5250] = 8'd142;
   assign soundFileAmplitudes [5251] = 8'd142;
   assign soundFileAmplitudes [5252] = 8'd140;
   assign soundFileAmplitudes [5253] = 8'd131;
   assign soundFileAmplitudes [5254] = 8'd128;
   assign soundFileAmplitudes [5255] = 8'd118;
   assign soundFileAmplitudes [5256] = 8'd124;
   assign soundFileAmplitudes [5257] = 8'd121;
   assign soundFileAmplitudes [5258] = 8'd123;
   assign soundFileAmplitudes [5259] = 8'd131;
   assign soundFileAmplitudes [5260] = 8'd124;
   assign soundFileAmplitudes [5261] = 8'd110;
   assign soundFileAmplitudes [5262] = 8'd99;
   assign soundFileAmplitudes [5263] = 8'd113;
   assign soundFileAmplitudes [5264] = 8'd120;
   assign soundFileAmplitudes [5265] = 8'd127;
   assign soundFileAmplitudes [5266] = 8'd136;
   assign soundFileAmplitudes [5267] = 8'd138;
   assign soundFileAmplitudes [5268] = 8'd140;
   assign soundFileAmplitudes [5269] = 8'd135;
   assign soundFileAmplitudes [5270] = 8'd142;
   assign soundFileAmplitudes [5271] = 8'd144;
   assign soundFileAmplitudes [5272] = 8'd145;
   assign soundFileAmplitudes [5273] = 8'd134;
   assign soundFileAmplitudes [5274] = 8'd121;
   assign soundFileAmplitudes [5275] = 8'd124;
   assign soundFileAmplitudes [5276] = 8'd106;
   assign soundFileAmplitudes [5277] = 8'd101;
   assign soundFileAmplitudes [5278] = 8'd103;
   assign soundFileAmplitudes [5279] = 8'd108;
   assign soundFileAmplitudes [5280] = 8'd114;
   assign soundFileAmplitudes [5281] = 8'd115;
   assign soundFileAmplitudes [5282] = 8'd121;
   assign soundFileAmplitudes [5283] = 8'd125;
   assign soundFileAmplitudes [5284] = 8'd123;
   assign soundFileAmplitudes [5285] = 8'd121;
   assign soundFileAmplitudes [5286] = 8'd125;
   assign soundFileAmplitudes [5287] = 8'd131;
   assign soundFileAmplitudes [5288] = 8'd126;
   assign soundFileAmplitudes [5289] = 8'd122;
   assign soundFileAmplitudes [5290] = 8'd127;
   assign soundFileAmplitudes [5291] = 8'd137;
   assign soundFileAmplitudes [5292] = 8'd138;
   assign soundFileAmplitudes [5293] = 8'd122;
   assign soundFileAmplitudes [5294] = 8'd124;
   assign soundFileAmplitudes [5295] = 8'd134;
   assign soundFileAmplitudes [5296] = 8'd129;
   assign soundFileAmplitudes [5297] = 8'd137;
   assign soundFileAmplitudes [5298] = 8'd142;
   assign soundFileAmplitudes [5299] = 8'd128;
   assign soundFileAmplitudes [5300] = 8'd125;
   assign soundFileAmplitudes [5301] = 8'd117;
   assign soundFileAmplitudes [5302] = 8'd125;
   assign soundFileAmplitudes [5303] = 8'd143;
   assign soundFileAmplitudes [5304] = 8'd149;
   assign soundFileAmplitudes [5305] = 8'd159;
   assign soundFileAmplitudes [5306] = 8'd158;
   assign soundFileAmplitudes [5307] = 8'd149;
   assign soundFileAmplitudes [5308] = 8'd145;
   assign soundFileAmplitudes [5309] = 8'd134;
   assign soundFileAmplitudes [5310] = 8'd132;
   assign soundFileAmplitudes [5311] = 8'd130;
   assign soundFileAmplitudes [5312] = 8'd110;
   assign soundFileAmplitudes [5313] = 8'd100;
   assign soundFileAmplitudes [5314] = 8'd92;
   assign soundFileAmplitudes [5315] = 8'd74;
   assign soundFileAmplitudes [5316] = 8'd68;
   assign soundFileAmplitudes [5317] = 8'd78;
   assign soundFileAmplitudes [5318] = 8'd96;
   assign soundFileAmplitudes [5319] = 8'd111;
   assign soundFileAmplitudes [5320] = 8'd115;
   assign soundFileAmplitudes [5321] = 8'd109;
   assign soundFileAmplitudes [5322] = 8'd108;
   assign soundFileAmplitudes [5323] = 8'd105;
   assign soundFileAmplitudes [5324] = 8'd113;
   assign soundFileAmplitudes [5325] = 8'd143;
   assign soundFileAmplitudes [5326] = 8'd160;
   assign soundFileAmplitudes [5327] = 8'd160;
   assign soundFileAmplitudes [5328] = 8'd153;
   assign soundFileAmplitudes [5329] = 8'd156;
   assign soundFileAmplitudes [5330] = 8'd178;
   assign soundFileAmplitudes [5331] = 8'd181;
   assign soundFileAmplitudes [5332] = 8'd157;
   assign soundFileAmplitudes [5333] = 8'd142;
   assign soundFileAmplitudes [5334] = 8'd131;
   assign soundFileAmplitudes [5335] = 8'd123;
   assign soundFileAmplitudes [5336] = 8'd127;
   assign soundFileAmplitudes [5337] = 8'd132;
   assign soundFileAmplitudes [5338] = 8'd135;
   assign soundFileAmplitudes [5339] = 8'd123;
   assign soundFileAmplitudes [5340] = 8'd111;
   assign soundFileAmplitudes [5341] = 8'd108;
   assign soundFileAmplitudes [5342] = 8'd123;
   assign soundFileAmplitudes [5343] = 8'd142;
   assign soundFileAmplitudes [5344] = 8'd145;
   assign soundFileAmplitudes [5345] = 8'd147;
   assign soundFileAmplitudes [5346] = 8'd139;
   assign soundFileAmplitudes [5347] = 8'd133;
   assign soundFileAmplitudes [5348] = 8'd122;
   assign soundFileAmplitudes [5349] = 8'd103;
   assign soundFileAmplitudes [5350] = 8'd99;
   assign soundFileAmplitudes [5351] = 8'd93;
   assign soundFileAmplitudes [5352] = 8'd91;
   assign soundFileAmplitudes [5353] = 8'd95;
   assign soundFileAmplitudes [5354] = 8'd86;
   assign soundFileAmplitudes [5355] = 8'd83;
   assign soundFileAmplitudes [5356] = 8'd80;
   assign soundFileAmplitudes [5357] = 8'd80;
   assign soundFileAmplitudes [5358] = 8'd100;
   assign soundFileAmplitudes [5359] = 8'd121;
   assign soundFileAmplitudes [5360] = 8'd145;
   assign soundFileAmplitudes [5361] = 8'd151;
   assign soundFileAmplitudes [5362] = 8'd150;
   assign soundFileAmplitudes [5363] = 8'd161;
   assign soundFileAmplitudes [5364] = 8'd173;
   assign soundFileAmplitudes [5365] = 8'd180;
   assign soundFileAmplitudes [5366] = 8'd162;
   assign soundFileAmplitudes [5367] = 8'd163;
   assign soundFileAmplitudes [5368] = 8'd161;
   assign soundFileAmplitudes [5369] = 8'd149;
   assign soundFileAmplitudes [5370] = 8'd133;
   assign soundFileAmplitudes [5371] = 8'd114;
   assign soundFileAmplitudes [5372] = 8'd113;
   assign soundFileAmplitudes [5373] = 8'd113;
   assign soundFileAmplitudes [5374] = 8'd121;
   assign soundFileAmplitudes [5375] = 8'd121;
   assign soundFileAmplitudes [5376] = 8'd115;
   assign soundFileAmplitudes [5377] = 8'd107;
   assign soundFileAmplitudes [5378] = 8'd102;
   assign soundFileAmplitudes [5379] = 8'd112;
   assign soundFileAmplitudes [5380] = 8'd122;
   assign soundFileAmplitudes [5381] = 8'd143;
   assign soundFileAmplitudes [5382] = 8'd147;
   assign soundFileAmplitudes [5383] = 8'd131;
   assign soundFileAmplitudes [5384] = 8'd128;
   assign soundFileAmplitudes [5385] = 8'd117;
   assign soundFileAmplitudes [5386] = 8'd120;
   assign soundFileAmplitudes [5387] = 8'd125;
   assign soundFileAmplitudes [5388] = 8'd101;
   assign soundFileAmplitudes [5389] = 8'd90;
   assign soundFileAmplitudes [5390] = 8'd83;
   assign soundFileAmplitudes [5391] = 8'd85;
   assign soundFileAmplitudes [5392] = 8'd92;
   assign soundFileAmplitudes [5393] = 8'd95;
   assign soundFileAmplitudes [5394] = 8'd111;
   assign soundFileAmplitudes [5395] = 8'd123;
   assign soundFileAmplitudes [5396] = 8'd137;
   assign soundFileAmplitudes [5397] = 8'd153;
   assign soundFileAmplitudes [5398] = 8'd152;
   assign soundFileAmplitudes [5399] = 8'd160;
   assign soundFileAmplitudes [5400] = 8'd163;
   assign soundFileAmplitudes [5401] = 8'd158;
   assign soundFileAmplitudes [5402] = 8'd161;
   assign soundFileAmplitudes [5403] = 8'd162;
   assign soundFileAmplitudes [5404] = 8'd157;
   assign soundFileAmplitudes [5405] = 8'd137;
   assign soundFileAmplitudes [5406] = 8'd129;
   assign soundFileAmplitudes [5407] = 8'd129;
   assign soundFileAmplitudes [5408] = 8'd128;
   assign soundFileAmplitudes [5409] = 8'd112;
   assign soundFileAmplitudes [5410] = 8'd99;
   assign soundFileAmplitudes [5411] = 8'd100;
   assign soundFileAmplitudes [5412] = 8'd101;
   assign soundFileAmplitudes [5413] = 8'd123;
   assign soundFileAmplitudes [5414] = 8'd123;
   assign soundFileAmplitudes [5415] = 8'd113;
   assign soundFileAmplitudes [5416] = 8'd114;
   assign soundFileAmplitudes [5417] = 8'd122;
   assign soundFileAmplitudes [5418] = 8'd121;
   assign soundFileAmplitudes [5419] = 8'd117;
   assign soundFileAmplitudes [5420] = 8'd128;
   assign soundFileAmplitudes [5421] = 8'd128;
   assign soundFileAmplitudes [5422] = 8'd122;
   assign soundFileAmplitudes [5423] = 8'd114;
   assign soundFileAmplitudes [5424] = 8'd103;
   assign soundFileAmplitudes [5425] = 8'd104;
   assign soundFileAmplitudes [5426] = 8'd106;
   assign soundFileAmplitudes [5427] = 8'd98;
   assign soundFileAmplitudes [5428] = 8'd104;
   assign soundFileAmplitudes [5429] = 8'd111;
   assign soundFileAmplitudes [5430] = 8'd123;
   assign soundFileAmplitudes [5431] = 8'd132;
   assign soundFileAmplitudes [5432] = 8'd135;
   assign soundFileAmplitudes [5433] = 8'd149;
   assign soundFileAmplitudes [5434] = 8'd156;
   assign soundFileAmplitudes [5435] = 8'd159;
   assign soundFileAmplitudes [5436] = 8'd164;
   assign soundFileAmplitudes [5437] = 8'd168;
   assign soundFileAmplitudes [5438] = 8'd168;
   assign soundFileAmplitudes [5439] = 8'd154;
   assign soundFileAmplitudes [5440] = 8'd129;
   assign soundFileAmplitudes [5441] = 8'd123;
   assign soundFileAmplitudes [5442] = 8'd127;
   assign soundFileAmplitudes [5443] = 8'd131;
   assign soundFileAmplitudes [5444] = 8'd121;
   assign soundFileAmplitudes [5445] = 8'd117;
   assign soundFileAmplitudes [5446] = 8'd121;
   assign soundFileAmplitudes [5447] = 8'd118;
   assign soundFileAmplitudes [5448] = 8'd124;
   assign soundFileAmplitudes [5449] = 8'd113;
   assign soundFileAmplitudes [5450] = 8'd100;
   assign soundFileAmplitudes [5451] = 8'd105;
   assign soundFileAmplitudes [5452] = 8'd115;
   assign soundFileAmplitudes [5453] = 8'd118;
   assign soundFileAmplitudes [5454] = 8'd118;
   assign soundFileAmplitudes [5455] = 8'd112;
   assign soundFileAmplitudes [5456] = 8'd107;
   assign soundFileAmplitudes [5457] = 8'd101;
   assign soundFileAmplitudes [5458] = 8'd110;
   assign soundFileAmplitudes [5459] = 8'd127;
   assign soundFileAmplitudes [5460] = 8'd141;
   assign soundFileAmplitudes [5461] = 8'd139;
   assign soundFileAmplitudes [5462] = 8'd123;
   assign soundFileAmplitudes [5463] = 8'd116;
   assign soundFileAmplitudes [5464] = 8'd119;
   assign soundFileAmplitudes [5465] = 8'd129;
   assign soundFileAmplitudes [5466] = 8'd136;
   assign soundFileAmplitudes [5467] = 8'd141;
   assign soundFileAmplitudes [5468] = 8'd139;
   assign soundFileAmplitudes [5469] = 8'd143;
   assign soundFileAmplitudes [5470] = 8'd151;
   assign soundFileAmplitudes [5471] = 8'd144;
   assign soundFileAmplitudes [5472] = 8'd136;
   assign soundFileAmplitudes [5473] = 8'd133;
   assign soundFileAmplitudes [5474] = 8'd129;
   assign soundFileAmplitudes [5475] = 8'd138;
   assign soundFileAmplitudes [5476] = 8'd147;
   assign soundFileAmplitudes [5477] = 8'd149;
   assign soundFileAmplitudes [5478] = 8'd153;
   assign soundFileAmplitudes [5479] = 8'd151;
   assign soundFileAmplitudes [5480] = 8'd135;
   assign soundFileAmplitudes [5481] = 8'd121;
   assign soundFileAmplitudes [5482] = 8'd115;
   assign soundFileAmplitudes [5483] = 8'd115;
   assign soundFileAmplitudes [5484] = 8'd120;
   assign soundFileAmplitudes [5485] = 8'd114;
   assign soundFileAmplitudes [5486] = 8'd112;
   assign soundFileAmplitudes [5487] = 8'd109;
   assign soundFileAmplitudes [5488] = 8'd112;
   assign soundFileAmplitudes [5489] = 8'd113;
   assign soundFileAmplitudes [5490] = 8'd96;
   assign soundFileAmplitudes [5491] = 8'd75;
   assign soundFileAmplitudes [5492] = 8'd73;
   assign soundFileAmplitudes [5493] = 8'd80;
   assign soundFileAmplitudes [5494] = 8'd93;
   assign soundFileAmplitudes [5495] = 8'd109;
   assign soundFileAmplitudes [5496] = 8'd124;
   assign soundFileAmplitudes [5497] = 8'd134;
   assign soundFileAmplitudes [5498] = 8'd135;
   assign soundFileAmplitudes [5499] = 8'd153;
   assign soundFileAmplitudes [5500] = 8'd178;
   assign soundFileAmplitudes [5501] = 8'd179;
   assign soundFileAmplitudes [5502] = 8'd167;
   assign soundFileAmplitudes [5503] = 8'd156;
   assign soundFileAmplitudes [5504] = 8'd156;
   assign soundFileAmplitudes [5505] = 8'd160;
   assign soundFileAmplitudes [5506] = 8'd150;
   assign soundFileAmplitudes [5507] = 8'd145;
   assign soundFileAmplitudes [5508] = 8'd138;
   assign soundFileAmplitudes [5509] = 8'd126;
   assign soundFileAmplitudes [5510] = 8'd114;
   assign soundFileAmplitudes [5511] = 8'd105;
   assign soundFileAmplitudes [5512] = 8'd104;
   assign soundFileAmplitudes [5513] = 8'd103;
   assign soundFileAmplitudes [5514] = 8'd100;
   assign soundFileAmplitudes [5515] = 8'd104;
   assign soundFileAmplitudes [5516] = 8'd112;
   assign soundFileAmplitudes [5517] = 8'd117;
   assign soundFileAmplitudes [5518] = 8'd123;
   assign soundFileAmplitudes [5519] = 8'd128;
   assign soundFileAmplitudes [5520] = 8'd128;
   assign soundFileAmplitudes [5521] = 8'd129;
   assign soundFileAmplitudes [5522] = 8'd120;
   assign soundFileAmplitudes [5523] = 8'd109;
   assign soundFileAmplitudes [5524] = 8'd113;
   assign soundFileAmplitudes [5525] = 8'd115;
   assign soundFileAmplitudes [5526] = 8'd103;
   assign soundFileAmplitudes [5527] = 8'd102;
   assign soundFileAmplitudes [5528] = 8'd123;
   assign soundFileAmplitudes [5529] = 8'd127;
   assign soundFileAmplitudes [5530] = 8'd109;
   assign soundFileAmplitudes [5531] = 8'd93;
   assign soundFileAmplitudes [5532] = 8'd97;
   assign soundFileAmplitudes [5533] = 8'd108;
   assign soundFileAmplitudes [5534] = 8'd136;
   assign soundFileAmplitudes [5535] = 8'd150;
   assign soundFileAmplitudes [5536] = 8'd151;
   assign soundFileAmplitudes [5537] = 8'd159;
   assign soundFileAmplitudes [5538] = 8'd159;
   assign soundFileAmplitudes [5539] = 8'd176;
   assign soundFileAmplitudes [5540] = 8'd185;
   assign soundFileAmplitudes [5541] = 8'd177;
   assign soundFileAmplitudes [5542] = 8'd157;
   assign soundFileAmplitudes [5543] = 8'd137;
   assign soundFileAmplitudes [5544] = 8'd121;
   assign soundFileAmplitudes [5545] = 8'd110;
   assign soundFileAmplitudes [5546] = 8'd98;
   assign soundFileAmplitudes [5547] = 8'd103;
   assign soundFileAmplitudes [5548] = 8'd106;
   assign soundFileAmplitudes [5549] = 8'd97;
   assign soundFileAmplitudes [5550] = 8'd94;
   assign soundFileAmplitudes [5551] = 8'd91;
   assign soundFileAmplitudes [5552] = 8'd96;
   assign soundFileAmplitudes [5553] = 8'd111;
   assign soundFileAmplitudes [5554] = 8'd122;
   assign soundFileAmplitudes [5555] = 8'd131;
   assign soundFileAmplitudes [5556] = 8'd136;
   assign soundFileAmplitudes [5557] = 8'd134;
   assign soundFileAmplitudes [5558] = 8'd139;
   assign soundFileAmplitudes [5559] = 8'd136;
   assign soundFileAmplitudes [5560] = 8'd134;
   assign soundFileAmplitudes [5561] = 8'd128;
   assign soundFileAmplitudes [5562] = 8'd125;
   assign soundFileAmplitudes [5563] = 8'd128;
   assign soundFileAmplitudes [5564] = 8'd125;
   assign soundFileAmplitudes [5565] = 8'd120;
   assign soundFileAmplitudes [5566] = 8'd110;
   assign soundFileAmplitudes [5567] = 8'd120;
   assign soundFileAmplitudes [5568] = 8'd124;
   assign soundFileAmplitudes [5569] = 8'd121;
   assign soundFileAmplitudes [5570] = 8'd119;
   assign soundFileAmplitudes [5571] = 8'd103;
   assign soundFileAmplitudes [5572] = 8'd96;
   assign soundFileAmplitudes [5573] = 8'd101;
   assign soundFileAmplitudes [5574] = 8'd116;
   assign soundFileAmplitudes [5575] = 8'd127;
   assign soundFileAmplitudes [5576] = 8'd134;
   assign soundFileAmplitudes [5577] = 8'd147;
   assign soundFileAmplitudes [5578] = 8'd152;
   assign soundFileAmplitudes [5579] = 8'd161;
   assign soundFileAmplitudes [5580] = 8'd161;
   assign soundFileAmplitudes [5581] = 8'd152;
   assign soundFileAmplitudes [5582] = 8'd147;
   assign soundFileAmplitudes [5583] = 8'd140;
   assign soundFileAmplitudes [5584] = 8'd139;
   assign soundFileAmplitudes [5585] = 8'd139;
   assign soundFileAmplitudes [5586] = 8'd128;
   assign soundFileAmplitudes [5587] = 8'd123;
   assign soundFileAmplitudes [5588] = 8'd127;
   assign soundFileAmplitudes [5589] = 8'd127;
   assign soundFileAmplitudes [5590] = 8'd122;
   assign soundFileAmplitudes [5591] = 8'd118;
   assign soundFileAmplitudes [5592] = 8'd110;
   assign soundFileAmplitudes [5593] = 8'd104;
   assign soundFileAmplitudes [5594] = 8'd104;
   assign soundFileAmplitudes [5595] = 8'd113;
   assign soundFileAmplitudes [5596] = 8'd123;
   assign soundFileAmplitudes [5597] = 8'd135;
   assign soundFileAmplitudes [5598] = 8'd137;
   assign soundFileAmplitudes [5599] = 8'd126;
   assign soundFileAmplitudes [5600] = 8'd122;
   assign soundFileAmplitudes [5601] = 8'd114;
   assign soundFileAmplitudes [5602] = 8'd106;
   assign soundFileAmplitudes [5603] = 8'd110;
   assign soundFileAmplitudes [5604] = 8'd122;
   assign soundFileAmplitudes [5605] = 8'd131;
   assign soundFileAmplitudes [5606] = 8'd136;
   assign soundFileAmplitudes [5607] = 8'd133;
   assign soundFileAmplitudes [5608] = 8'd132;
   assign soundFileAmplitudes [5609] = 8'd125;
   assign soundFileAmplitudes [5610] = 8'd128;
   assign soundFileAmplitudes [5611] = 8'd125;
   assign soundFileAmplitudes [5612] = 8'd109;
   assign soundFileAmplitudes [5613] = 8'd111;
   assign soundFileAmplitudes [5614] = 8'd112;
   assign soundFileAmplitudes [5615] = 8'd118;
   assign soundFileAmplitudes [5616] = 8'd130;
   assign soundFileAmplitudes [5617] = 8'd136;
   assign soundFileAmplitudes [5618] = 8'd147;
   assign soundFileAmplitudes [5619] = 8'd156;
   assign soundFileAmplitudes [5620] = 8'd154;
   assign soundFileAmplitudes [5621] = 8'd150;
   assign soundFileAmplitudes [5622] = 8'd135;
   assign soundFileAmplitudes [5623] = 8'd125;
   assign soundFileAmplitudes [5624] = 8'd129;
   assign soundFileAmplitudes [5625] = 8'd131;
   assign soundFileAmplitudes [5626] = 8'd133;
   assign soundFileAmplitudes [5627] = 8'd134;
   assign soundFileAmplitudes [5628] = 8'd122;
   assign soundFileAmplitudes [5629] = 8'd114;
   assign soundFileAmplitudes [5630] = 8'd112;
   assign soundFileAmplitudes [5631] = 8'd110;
   assign soundFileAmplitudes [5632] = 8'd116;
   assign soundFileAmplitudes [5633] = 8'd115;
   assign soundFileAmplitudes [5634] = 8'd125;
   assign soundFileAmplitudes [5635] = 8'd126;
   assign soundFileAmplitudes [5636] = 8'd130;
   assign soundFileAmplitudes [5637] = 8'd134;
   assign soundFileAmplitudes [5638] = 8'd123;
   assign soundFileAmplitudes [5639] = 8'd129;
   assign soundFileAmplitudes [5640] = 8'd140;
   assign soundFileAmplitudes [5641] = 8'd140;
   assign soundFileAmplitudes [5642] = 8'd134;
   assign soundFileAmplitudes [5643] = 8'd133;
   assign soundFileAmplitudes [5644] = 8'd132;
   assign soundFileAmplitudes [5645] = 8'd138;
   assign soundFileAmplitudes [5646] = 8'd128;
   assign soundFileAmplitudes [5647] = 8'd117;
   assign soundFileAmplitudes [5648] = 8'd117;
   assign soundFileAmplitudes [5649] = 8'd116;
   assign soundFileAmplitudes [5650] = 8'd121;
   assign soundFileAmplitudes [5651] = 8'd110;
   assign soundFileAmplitudes [5652] = 8'd109;
   assign soundFileAmplitudes [5653] = 8'd112;
   assign soundFileAmplitudes [5654] = 8'd106;
   assign soundFileAmplitudes [5655] = 8'd97;
   assign soundFileAmplitudes [5656] = 8'd96;
   assign soundFileAmplitudes [5657] = 8'd102;
   assign soundFileAmplitudes [5658] = 8'd112;
   assign soundFileAmplitudes [5659] = 8'd119;
   assign soundFileAmplitudes [5660] = 8'd125;
   assign soundFileAmplitudes [5661] = 8'd138;
   assign soundFileAmplitudes [5662] = 8'd142;
   assign soundFileAmplitudes [5663] = 8'd137;
   assign soundFileAmplitudes [5664] = 8'd131;
   assign soundFileAmplitudes [5665] = 8'd126;
   assign soundFileAmplitudes [5666] = 8'd127;
   assign soundFileAmplitudes [5667] = 8'd119;
   assign soundFileAmplitudes [5668] = 8'd125;
   assign soundFileAmplitudes [5669] = 8'd140;
   assign soundFileAmplitudes [5670] = 8'd145;
   assign soundFileAmplitudes [5671] = 8'd150;
   assign soundFileAmplitudes [5672] = 8'd131;
   assign soundFileAmplitudes [5673] = 8'd126;
   assign soundFileAmplitudes [5674] = 8'd124;
   assign soundFileAmplitudes [5675] = 8'd124;
   assign soundFileAmplitudes [5676] = 8'd130;
   assign soundFileAmplitudes [5677] = 8'd134;
   assign soundFileAmplitudes [5678] = 8'd139;
   assign soundFileAmplitudes [5679] = 8'd141;
   assign soundFileAmplitudes [5680] = 8'd137;
   assign soundFileAmplitudes [5681] = 8'd133;
   assign soundFileAmplitudes [5682] = 8'd133;
   assign soundFileAmplitudes [5683] = 8'd132;
   assign soundFileAmplitudes [5684] = 8'd132;
   assign soundFileAmplitudes [5685] = 8'd129;
   assign soundFileAmplitudes [5686] = 8'd119;
   assign soundFileAmplitudes [5687] = 8'd112;
   assign soundFileAmplitudes [5688] = 8'd116;
   assign soundFileAmplitudes [5689] = 8'd123;
   assign soundFileAmplitudes [5690] = 8'd134;
   assign soundFileAmplitudes [5691] = 8'd129;
   assign soundFileAmplitudes [5692] = 8'd115;
   assign soundFileAmplitudes [5693] = 8'd105;
   assign soundFileAmplitudes [5694] = 8'd103;
   assign soundFileAmplitudes [5695] = 8'd102;
   assign soundFileAmplitudes [5696] = 8'd97;
   assign soundFileAmplitudes [5697] = 8'd99;
   assign soundFileAmplitudes [5698] = 8'd112;
   assign soundFileAmplitudes [5699] = 8'd117;
   assign soundFileAmplitudes [5700] = 8'd118;
   assign soundFileAmplitudes [5701] = 8'd116;
   assign soundFileAmplitudes [5702] = 8'd117;
   assign soundFileAmplitudes [5703] = 8'd125;
   assign soundFileAmplitudes [5704] = 8'd137;
   assign soundFileAmplitudes [5705] = 8'd147;
   assign soundFileAmplitudes [5706] = 8'd146;
   assign soundFileAmplitudes [5707] = 8'd138;
   assign soundFileAmplitudes [5708] = 8'd129;
   assign soundFileAmplitudes [5709] = 8'd118;
   assign soundFileAmplitudes [5710] = 8'd116;
   assign soundFileAmplitudes [5711] = 8'd132;
   assign soundFileAmplitudes [5712] = 8'd132;
   assign soundFileAmplitudes [5713] = 8'd133;
   assign soundFileAmplitudes [5714] = 8'd131;
   assign soundFileAmplitudes [5715] = 8'd126;
   assign soundFileAmplitudes [5716] = 8'd127;
   assign soundFileAmplitudes [5717] = 8'd136;
   assign soundFileAmplitudes [5718] = 8'd133;
   assign soundFileAmplitudes [5719] = 8'd136;
   assign soundFileAmplitudes [5720] = 8'd138;
   assign soundFileAmplitudes [5721] = 8'd132;
   assign soundFileAmplitudes [5722] = 8'd137;
   assign soundFileAmplitudes [5723] = 8'd144;
   assign soundFileAmplitudes [5724] = 8'd152;
   assign soundFileAmplitudes [5725] = 8'd147;
   assign soundFileAmplitudes [5726] = 8'd151;
   assign soundFileAmplitudes [5727] = 8'd142;
   assign soundFileAmplitudes [5728] = 8'd133;
   assign soundFileAmplitudes [5729] = 8'd122;
   assign soundFileAmplitudes [5730] = 8'd117;
   assign soundFileAmplitudes [5731] = 8'd114;
   assign soundFileAmplitudes [5732] = 8'd115;
   assign soundFileAmplitudes [5733] = 8'd120;
   assign soundFileAmplitudes [5734] = 8'd116;
   assign soundFileAmplitudes [5735] = 8'd111;
   assign soundFileAmplitudes [5736] = 8'd111;
   assign soundFileAmplitudes [5737] = 8'd121;
   assign soundFileAmplitudes [5738] = 8'd127;
   assign soundFileAmplitudes [5739] = 8'd125;
   assign soundFileAmplitudes [5740] = 8'd114;
   assign soundFileAmplitudes [5741] = 8'd102;
   assign soundFileAmplitudes [5742] = 8'd96;
   assign soundFileAmplitudes [5743] = 8'd109;
   assign soundFileAmplitudes [5744] = 8'd111;
   assign soundFileAmplitudes [5745] = 8'd110;
   assign soundFileAmplitudes [5746] = 8'd114;
   assign soundFileAmplitudes [5747] = 8'd115;
   assign soundFileAmplitudes [5748] = 8'd131;
   assign soundFileAmplitudes [5749] = 8'd145;
   assign soundFileAmplitudes [5750] = 8'd144;
   assign soundFileAmplitudes [5751] = 8'd139;
   assign soundFileAmplitudes [5752] = 8'd136;
   assign soundFileAmplitudes [5753] = 8'd143;
   assign soundFileAmplitudes [5754] = 8'd148;
   assign soundFileAmplitudes [5755] = 8'd149;
   assign soundFileAmplitudes [5756] = 8'd150;
   assign soundFileAmplitudes [5757] = 8'd150;
   assign soundFileAmplitudes [5758] = 8'd148;
   assign soundFileAmplitudes [5759] = 8'd134;
   assign soundFileAmplitudes [5760] = 8'd126;
   assign soundFileAmplitudes [5761] = 8'd124;
   assign soundFileAmplitudes [5762] = 8'd126;
   assign soundFileAmplitudes [5763] = 8'd125;
   assign soundFileAmplitudes [5764] = 8'd117;
   assign soundFileAmplitudes [5765] = 8'd122;
   assign soundFileAmplitudes [5766] = 8'd120;
   assign soundFileAmplitudes [5767] = 8'd128;
   assign soundFileAmplitudes [5768] = 8'd131;
   assign soundFileAmplitudes [5769] = 8'd131;
   assign soundFileAmplitudes [5770] = 8'd127;
   assign soundFileAmplitudes [5771] = 8'd118;
   assign soundFileAmplitudes [5772] = 8'd123;
   assign soundFileAmplitudes [5773] = 8'd123;
   assign soundFileAmplitudes [5774] = 8'd121;
   assign soundFileAmplitudes [5775] = 8'd117;
   assign soundFileAmplitudes [5776] = 8'd121;
   assign soundFileAmplitudes [5777] = 8'd119;
   assign soundFileAmplitudes [5778] = 8'd116;
   assign soundFileAmplitudes [5779] = 8'd108;
   assign soundFileAmplitudes [5780] = 8'd95;
   assign soundFileAmplitudes [5781] = 8'd88;
   assign soundFileAmplitudes [5782] = 8'd96;
   assign soundFileAmplitudes [5783] = 8'd116;
   assign soundFileAmplitudes [5784] = 8'd128;
   assign soundFileAmplitudes [5785] = 8'd132;
   assign soundFileAmplitudes [5786] = 8'd139;
   assign soundFileAmplitudes [5787] = 8'd128;
   assign soundFileAmplitudes [5788] = 8'd131;
   assign soundFileAmplitudes [5789] = 8'd143;
   assign soundFileAmplitudes [5790] = 8'd139;
   assign soundFileAmplitudes [5791] = 8'd141;
   assign soundFileAmplitudes [5792] = 8'd134;
   assign soundFileAmplitudes [5793] = 8'd137;
   assign soundFileAmplitudes [5794] = 8'd140;
   assign soundFileAmplitudes [5795] = 8'd130;
   assign soundFileAmplitudes [5796] = 8'd119;
   assign soundFileAmplitudes [5797] = 8'd125;
   assign soundFileAmplitudes [5798] = 8'd129;
   assign soundFileAmplitudes [5799] = 8'd124;
   assign soundFileAmplitudes [5800] = 8'd117;
   assign soundFileAmplitudes [5801] = 8'd113;
   assign soundFileAmplitudes [5802] = 8'd128;
   assign soundFileAmplitudes [5803] = 8'd136;
   assign soundFileAmplitudes [5804] = 8'd143;
   assign soundFileAmplitudes [5805] = 8'd147;
   assign soundFileAmplitudes [5806] = 8'd142;
   assign soundFileAmplitudes [5807] = 8'd140;
   assign soundFileAmplitudes [5808] = 8'd133;
   assign soundFileAmplitudes [5809] = 8'd132;
   assign soundFileAmplitudes [5810] = 8'd122;
   assign soundFileAmplitudes [5811] = 8'd115;
   assign soundFileAmplitudes [5812] = 8'd116;
   assign soundFileAmplitudes [5813] = 8'd108;
   assign soundFileAmplitudes [5814] = 8'd103;
   assign soundFileAmplitudes [5815] = 8'd98;
   assign soundFileAmplitudes [5816] = 8'd102;
   assign soundFileAmplitudes [5817] = 8'd104;
   assign soundFileAmplitudes [5818] = 8'd110;
   assign soundFileAmplitudes [5819] = 8'd107;
   assign soundFileAmplitudes [5820] = 8'd109;
   assign soundFileAmplitudes [5821] = 8'd128;
   assign soundFileAmplitudes [5822] = 8'd136;
   assign soundFileAmplitudes [5823] = 8'd140;
   assign soundFileAmplitudes [5824] = 8'd140;
   assign soundFileAmplitudes [5825] = 8'd139;
   assign soundFileAmplitudes [5826] = 8'd143;
   assign soundFileAmplitudes [5827] = 8'd148;
   assign soundFileAmplitudes [5828] = 8'd148;
   assign soundFileAmplitudes [5829] = 8'd140;
   assign soundFileAmplitudes [5830] = 8'd131;
   assign soundFileAmplitudes [5831] = 8'd117;
   assign soundFileAmplitudes [5832] = 8'd114;
   assign soundFileAmplitudes [5833] = 8'd115;
   assign soundFileAmplitudes [5834] = 8'd116;
   assign soundFileAmplitudes [5835] = 8'd117;
   assign soundFileAmplitudes [5836] = 8'd112;
   assign soundFileAmplitudes [5837] = 8'd120;
   assign soundFileAmplitudes [5838] = 8'd117;
   assign soundFileAmplitudes [5839] = 8'd118;
   assign soundFileAmplitudes [5840] = 8'd124;
   assign soundFileAmplitudes [5841] = 8'd134;
   assign soundFileAmplitudes [5842] = 8'd144;
   assign soundFileAmplitudes [5843] = 8'd150;
   assign soundFileAmplitudes [5844] = 8'd150;
   assign soundFileAmplitudes [5845] = 8'd150;
   assign soundFileAmplitudes [5846] = 8'd139;
   assign soundFileAmplitudes [5847] = 8'd129;
   assign soundFileAmplitudes [5848] = 8'd127;
   assign soundFileAmplitudes [5849] = 8'd131;
   assign soundFileAmplitudes [5850] = 8'd137;
   assign soundFileAmplitudes [5851] = 8'd121;
   assign soundFileAmplitudes [5852] = 8'd118;
   assign soundFileAmplitudes [5853] = 8'd105;
   assign soundFileAmplitudes [5854] = 8'd106;
   assign soundFileAmplitudes [5855] = 8'd121;
   assign soundFileAmplitudes [5856] = 8'd124;
   assign soundFileAmplitudes [5857] = 8'd128;
   assign soundFileAmplitudes [5858] = 8'd107;
   assign soundFileAmplitudes [5859] = 8'd90;
   assign soundFileAmplitudes [5860] = 8'd101;
   assign soundFileAmplitudes [5861] = 8'd126;
   assign soundFileAmplitudes [5862] = 8'd132;
   assign soundFileAmplitudes [5863] = 8'd129;
   assign soundFileAmplitudes [5864] = 8'd131;
   assign soundFileAmplitudes [5865] = 8'd131;
   assign soundFileAmplitudes [5866] = 8'd131;
   assign soundFileAmplitudes [5867] = 8'd132;
   assign soundFileAmplitudes [5868] = 8'd132;
   assign soundFileAmplitudes [5869] = 8'd129;
   assign soundFileAmplitudes [5870] = 8'd119;
   assign soundFileAmplitudes [5871] = 8'd126;
   assign soundFileAmplitudes [5872] = 8'd136;
   assign soundFileAmplitudes [5873] = 8'd141;
   assign soundFileAmplitudes [5874] = 8'd140;
   assign soundFileAmplitudes [5875] = 8'd131;
   assign soundFileAmplitudes [5876] = 8'd130;
   assign soundFileAmplitudes [5877] = 8'd129;
   assign soundFileAmplitudes [5878] = 8'd128;
   assign soundFileAmplitudes [5879] = 8'd123;
   assign soundFileAmplitudes [5880] = 8'd130;
   assign soundFileAmplitudes [5881] = 8'd135;
   assign soundFileAmplitudes [5882] = 8'd146;
   assign soundFileAmplitudes [5883] = 8'd139;
   assign soundFileAmplitudes [5884] = 8'd135;
   assign soundFileAmplitudes [5885] = 8'd130;
   assign soundFileAmplitudes [5886] = 8'd128;
   assign soundFileAmplitudes [5887] = 8'd128;
   assign soundFileAmplitudes [5888] = 8'd125;
   assign soundFileAmplitudes [5889] = 8'd123;
   assign soundFileAmplitudes [5890] = 8'd112;
   assign soundFileAmplitudes [5891] = 8'd121;
   assign soundFileAmplitudes [5892] = 8'd123;
   assign soundFileAmplitudes [5893] = 8'd133;
   assign soundFileAmplitudes [5894] = 8'd119;
   assign soundFileAmplitudes [5895] = 8'd95;
   assign soundFileAmplitudes [5896] = 8'd94;
   assign soundFileAmplitudes [5897] = 8'd111;
   assign soundFileAmplitudes [5898] = 8'd114;
   assign soundFileAmplitudes [5899] = 8'd110;
   assign soundFileAmplitudes [5900] = 8'd117;
   assign soundFileAmplitudes [5901] = 8'd118;
   assign soundFileAmplitudes [5902] = 8'd130;
   assign soundFileAmplitudes [5903] = 8'd143;
   assign soundFileAmplitudes [5904] = 8'd148;
   assign soundFileAmplitudes [5905] = 8'd144;
   assign soundFileAmplitudes [5906] = 8'd136;
   assign soundFileAmplitudes [5907] = 8'd130;
   assign soundFileAmplitudes [5908] = 8'd130;
   assign soundFileAmplitudes [5909] = 8'd141;
   assign soundFileAmplitudes [5910] = 8'd144;
   assign soundFileAmplitudes [5911] = 8'd136;
   assign soundFileAmplitudes [5912] = 8'd129;
   assign soundFileAmplitudes [5913] = 8'd128;
   assign soundFileAmplitudes [5914] = 8'd133;
   assign soundFileAmplitudes [5915] = 8'd127;
   assign soundFileAmplitudes [5916] = 8'd123;
   assign soundFileAmplitudes [5917] = 8'd115;
   assign soundFileAmplitudes [5918] = 8'd121;
   assign soundFileAmplitudes [5919] = 8'd126;
   assign soundFileAmplitudes [5920] = 8'd133;
   assign soundFileAmplitudes [5921] = 8'd137;
   assign soundFileAmplitudes [5922] = 8'd135;
   assign soundFileAmplitudes [5923] = 8'd127;
   assign soundFileAmplitudes [5924] = 8'd113;
   assign soundFileAmplitudes [5925] = 8'd107;
   assign soundFileAmplitudes [5926] = 8'd117;
   assign soundFileAmplitudes [5927] = 8'd129;
   assign soundFileAmplitudes [5928] = 8'd110;
   assign soundFileAmplitudes [5929] = 8'd119;
   assign soundFileAmplitudes [5930] = 8'd115;
   assign soundFileAmplitudes [5931] = 8'd113;
   assign soundFileAmplitudes [5932] = 8'd110;
   assign soundFileAmplitudes [5933] = 8'd88;
   assign soundFileAmplitudes [5934] = 8'd97;
   assign soundFileAmplitudes [5935] = 8'd114;
   assign soundFileAmplitudes [5936] = 8'd122;
   assign soundFileAmplitudes [5937] = 8'd125;
   assign soundFileAmplitudes [5938] = 8'd130;
   assign soundFileAmplitudes [5939] = 8'd122;
   assign soundFileAmplitudes [5940] = 8'd128;
   assign soundFileAmplitudes [5941] = 8'd141;
   assign soundFileAmplitudes [5942] = 8'd151;
   assign soundFileAmplitudes [5943] = 8'd159;
   assign soundFileAmplitudes [5944] = 8'd151;
   assign soundFileAmplitudes [5945] = 8'd136;
   assign soundFileAmplitudes [5946] = 8'd130;
   assign soundFileAmplitudes [5947] = 8'd134;
   assign soundFileAmplitudes [5948] = 8'd135;
   assign soundFileAmplitudes [5949] = 8'd139;
   assign soundFileAmplitudes [5950] = 8'd141;
   assign soundFileAmplitudes [5951] = 8'd132;
   assign soundFileAmplitudes [5952] = 8'd122;
   assign soundFileAmplitudes [5953] = 8'd114;
   assign soundFileAmplitudes [5954] = 8'd111;
   assign soundFileAmplitudes [5955] = 8'd115;
   assign soundFileAmplitudes [5956] = 8'd115;
   assign soundFileAmplitudes [5957] = 8'd126;
   assign soundFileAmplitudes [5958] = 8'd139;
   assign soundFileAmplitudes [5959] = 8'd131;
   assign soundFileAmplitudes [5960] = 8'd117;
   assign soundFileAmplitudes [5961] = 8'd117;
   assign soundFileAmplitudes [5962] = 8'd113;
   assign soundFileAmplitudes [5963] = 8'd123;
   assign soundFileAmplitudes [5964] = 8'd130;
   assign soundFileAmplitudes [5965] = 8'd120;
   assign soundFileAmplitudes [5966] = 8'd133;
   assign soundFileAmplitudes [5967] = 8'd134;
   assign soundFileAmplitudes [5968] = 8'd134;
   assign soundFileAmplitudes [5969] = 8'd125;
   assign soundFileAmplitudes [5970] = 8'd101;
   assign soundFileAmplitudes [5971] = 8'd107;
   assign soundFileAmplitudes [5972] = 8'd115;
   assign soundFileAmplitudes [5973] = 8'd130;
   assign soundFileAmplitudes [5974] = 8'd134;
   assign soundFileAmplitudes [5975] = 8'd111;
   assign soundFileAmplitudes [5976] = 8'd99;
   assign soundFileAmplitudes [5977] = 8'd99;
   assign soundFileAmplitudes [5978] = 8'd107;
   assign soundFileAmplitudes [5979] = 8'd133;
   assign soundFileAmplitudes [5980] = 8'd150;
   assign soundFileAmplitudes [5981] = 8'd143;
   assign soundFileAmplitudes [5982] = 8'd130;
   assign soundFileAmplitudes [5983] = 8'd131;
   assign soundFileAmplitudes [5984] = 8'd139;
   assign soundFileAmplitudes [5985] = 8'd150;
   assign soundFileAmplitudes [5986] = 8'd151;
   assign soundFileAmplitudes [5987] = 8'd147;
   assign soundFileAmplitudes [5988] = 8'd145;
   assign soundFileAmplitudes [5989] = 8'd138;
   assign soundFileAmplitudes [5990] = 8'd131;
   assign soundFileAmplitudes [5991] = 8'd115;
   assign soundFileAmplitudes [5992] = 8'd112;
   assign soundFileAmplitudes [5993] = 8'd126;
   assign soundFileAmplitudes [5994] = 8'd132;
   assign soundFileAmplitudes [5995] = 8'd124;
   assign soundFileAmplitudes [5996] = 8'd118;
   assign soundFileAmplitudes [5997] = 8'd104;
   assign soundFileAmplitudes [5998] = 8'd103;
   assign soundFileAmplitudes [5999] = 8'd113;
   assign soundFileAmplitudes [6000] = 8'd134;
   assign soundFileAmplitudes [6001] = 8'd137;
   assign soundFileAmplitudes [6002] = 8'd122;
   assign soundFileAmplitudes [6003] = 8'd134;
   assign soundFileAmplitudes [6004] = 8'd131;
   assign soundFileAmplitudes [6005] = 8'd144;
   assign soundFileAmplitudes [6006] = 8'd131;
   assign soundFileAmplitudes [6007] = 8'd114;
   assign soundFileAmplitudes [6008] = 8'd123;
   assign soundFileAmplitudes [6009] = 8'd118;
   assign soundFileAmplitudes [6010] = 8'd123;
   assign soundFileAmplitudes [6011] = 8'd110;
   assign soundFileAmplitudes [6012] = 8'd104;
   assign soundFileAmplitudes [6013] = 8'd107;
   assign soundFileAmplitudes [6014] = 8'd112;
   assign soundFileAmplitudes [6015] = 8'd134;
   assign soundFileAmplitudes [6016] = 8'd146;
   assign soundFileAmplitudes [6017] = 8'd150;
   assign soundFileAmplitudes [6018] = 8'd149;
   assign soundFileAmplitudes [6019] = 8'd141;
   assign soundFileAmplitudes [6020] = 8'd147;
   assign soundFileAmplitudes [6021] = 8'd146;
   assign soundFileAmplitudes [6022] = 8'd143;
   assign soundFileAmplitudes [6023] = 8'd143;
   assign soundFileAmplitudes [6024] = 8'd133;
   assign soundFileAmplitudes [6025] = 8'd135;
   assign soundFileAmplitudes [6026] = 8'd130;
   assign soundFileAmplitudes [6027] = 8'd123;
   assign soundFileAmplitudes [6028] = 8'd117;
   assign soundFileAmplitudes [6029] = 8'd107;
   assign soundFileAmplitudes [6030] = 8'd106;
   assign soundFileAmplitudes [6031] = 8'd107;
   assign soundFileAmplitudes [6032] = 8'd116;
   assign soundFileAmplitudes [6033] = 8'd116;
   assign soundFileAmplitudes [6034] = 8'd109;
   assign soundFileAmplitudes [6035] = 8'd111;
   assign soundFileAmplitudes [6036] = 8'd123;
   assign soundFileAmplitudes [6037] = 8'd129;
   assign soundFileAmplitudes [6038] = 8'd135;
   assign soundFileAmplitudes [6039] = 8'd133;
   assign soundFileAmplitudes [6040] = 8'd128;
   assign soundFileAmplitudes [6041] = 8'd140;
   assign soundFileAmplitudes [6042] = 8'd138;
   assign soundFileAmplitudes [6043] = 8'd132;
   assign soundFileAmplitudes [6044] = 8'd123;
   assign soundFileAmplitudes [6045] = 8'd107;
   assign soundFileAmplitudes [6046] = 8'd107;
   assign soundFileAmplitudes [6047] = 8'd116;
   assign soundFileAmplitudes [6048] = 8'd111;
   assign soundFileAmplitudes [6049] = 8'd110;
   assign soundFileAmplitudes [6050] = 8'd111;
   assign soundFileAmplitudes [6051] = 8'd107;
   assign soundFileAmplitudes [6052] = 8'd122;
   assign soundFileAmplitudes [6053] = 8'd141;
   assign soundFileAmplitudes [6054] = 8'd147;
   assign soundFileAmplitudes [6055] = 8'd147;
   assign soundFileAmplitudes [6056] = 8'd142;
   assign soundFileAmplitudes [6057] = 8'd136;
   assign soundFileAmplitudes [6058] = 8'd146;
   assign soundFileAmplitudes [6059] = 8'd153;
   assign soundFileAmplitudes [6060] = 8'd150;
   assign soundFileAmplitudes [6061] = 8'd139;
   assign soundFileAmplitudes [6062] = 8'd137;
   assign soundFileAmplitudes [6063] = 8'd127;
   assign soundFileAmplitudes [6064] = 8'd110;
   assign soundFileAmplitudes [6065] = 8'd111;
   assign soundFileAmplitudes [6066] = 8'd105;
   assign soundFileAmplitudes [6067] = 8'd101;
   assign soundFileAmplitudes [6068] = 8'd111;
   assign soundFileAmplitudes [6069] = 8'd118;
   assign soundFileAmplitudes [6070] = 8'd116;
   assign soundFileAmplitudes [6071] = 8'd118;
   assign soundFileAmplitudes [6072] = 8'd128;
   assign soundFileAmplitudes [6073] = 8'd132;
   assign soundFileAmplitudes [6074] = 8'd136;
   assign soundFileAmplitudes [6075] = 8'd143;
   assign soundFileAmplitudes [6076] = 8'd130;
   assign soundFileAmplitudes [6077] = 8'd134;
   assign soundFileAmplitudes [6078] = 8'd143;
   assign soundFileAmplitudes [6079] = 8'd133;
   assign soundFileAmplitudes [6080] = 8'd134;
   assign soundFileAmplitudes [6081] = 8'd125;
   assign soundFileAmplitudes [6082] = 8'd110;
   assign soundFileAmplitudes [6083] = 8'd106;
   assign soundFileAmplitudes [6084] = 8'd99;
   assign soundFileAmplitudes [6085] = 8'd99;
   assign soundFileAmplitudes [6086] = 8'd103;
   assign soundFileAmplitudes [6087] = 8'd112;
   assign soundFileAmplitudes [6088] = 8'd114;
   assign soundFileAmplitudes [6089] = 8'd122;
   assign soundFileAmplitudes [6090] = 8'd131;
   assign soundFileAmplitudes [6091] = 8'd131;
   assign soundFileAmplitudes [6092] = 8'd143;
   assign soundFileAmplitudes [6093] = 8'd138;
   assign soundFileAmplitudes [6094] = 8'd137;
   assign soundFileAmplitudes [6095] = 8'd143;
   assign soundFileAmplitudes [6096] = 8'd148;
   assign soundFileAmplitudes [6097] = 8'd151;
   assign soundFileAmplitudes [6098] = 8'd149;
   assign soundFileAmplitudes [6099] = 8'd141;
   assign soundFileAmplitudes [6100] = 8'd118;
   assign soundFileAmplitudes [6101] = 8'd113;
   assign soundFileAmplitudes [6102] = 8'd106;
   assign soundFileAmplitudes [6103] = 8'd98;
   assign soundFileAmplitudes [6104] = 8'd98;
   assign soundFileAmplitudes [6105] = 8'd98;
   assign soundFileAmplitudes [6106] = 8'd110;
   assign soundFileAmplitudes [6107] = 8'd123;
   assign soundFileAmplitudes [6108] = 8'd123;
   assign soundFileAmplitudes [6109] = 8'd128;
   assign soundFileAmplitudes [6110] = 8'd132;
   assign soundFileAmplitudes [6111] = 8'd132;
   assign soundFileAmplitudes [6112] = 8'd135;
   assign soundFileAmplitudes [6113] = 8'd144;
   assign soundFileAmplitudes [6114] = 8'd146;
   assign soundFileAmplitudes [6115] = 8'd135;
   assign soundFileAmplitudes [6116] = 8'd131;
   assign soundFileAmplitudes [6117] = 8'd139;
   assign soundFileAmplitudes [6118] = 8'd144;
   assign soundFileAmplitudes [6119] = 8'd132;
   assign soundFileAmplitudes [6120] = 8'd109;
   assign soundFileAmplitudes [6121] = 8'd96;
   assign soundFileAmplitudes [6122] = 8'd107;
   assign soundFileAmplitudes [6123] = 8'd120;
   assign soundFileAmplitudes [6124] = 8'd125;
   assign soundFileAmplitudes [6125] = 8'd118;
   assign soundFileAmplitudes [6126] = 8'd118;
   assign soundFileAmplitudes [6127] = 8'd125;
   assign soundFileAmplitudes [6128] = 8'd142;
   assign soundFileAmplitudes [6129] = 8'd156;
   assign soundFileAmplitudes [6130] = 8'd159;
   assign soundFileAmplitudes [6131] = 8'd159;
   assign soundFileAmplitudes [6132] = 8'd151;
   assign soundFileAmplitudes [6133] = 8'd151;
   assign soundFileAmplitudes [6134] = 8'd141;
   assign soundFileAmplitudes [6135] = 8'd141;
   assign soundFileAmplitudes [6136] = 8'd133;
   assign soundFileAmplitudes [6137] = 8'd120;
   assign soundFileAmplitudes [6138] = 8'd120;
   assign soundFileAmplitudes [6139] = 8'd107;
   assign soundFileAmplitudes [6140] = 8'd92;
   assign soundFileAmplitudes [6141] = 8'd87;
   assign soundFileAmplitudes [6142] = 8'd102;
   assign soundFileAmplitudes [6143] = 8'd121;
   assign soundFileAmplitudes [6144] = 8'd119;
   assign soundFileAmplitudes [6145] = 8'd113;
   assign soundFileAmplitudes [6146] = 8'd116;
   assign soundFileAmplitudes [6147] = 8'd119;
   assign soundFileAmplitudes [6148] = 8'd114;
   assign soundFileAmplitudes [6149] = 8'd120;
   assign soundFileAmplitudes [6150] = 8'd129;
   assign soundFileAmplitudes [6151] = 8'd132;
   assign soundFileAmplitudes [6152] = 8'd140;
   assign soundFileAmplitudes [6153] = 8'd134;
   assign soundFileAmplitudes [6154] = 8'd135;
   assign soundFileAmplitudes [6155] = 8'd130;
   assign soundFileAmplitudes [6156] = 8'd120;
   assign soundFileAmplitudes [6157] = 8'd119;
   assign soundFileAmplitudes [6158] = 8'd103;
   assign soundFileAmplitudes [6159] = 8'd103;
   assign soundFileAmplitudes [6160] = 8'd117;
   assign soundFileAmplitudes [6161] = 8'd119;
   assign soundFileAmplitudes [6162] = 8'd113;
   assign soundFileAmplitudes [6163] = 8'd120;
   assign soundFileAmplitudes [6164] = 8'd136;
   assign soundFileAmplitudes [6165] = 8'd151;
   assign soundFileAmplitudes [6166] = 8'd157;
   assign soundFileAmplitudes [6167] = 8'd156;
   assign soundFileAmplitudes [6168] = 8'd152;
   assign soundFileAmplitudes [6169] = 8'd145;
   assign soundFileAmplitudes [6170] = 8'd143;
   assign soundFileAmplitudes [6171] = 8'd142;
   assign soundFileAmplitudes [6172] = 8'd146;
   assign soundFileAmplitudes [6173] = 8'd138;
   assign soundFileAmplitudes [6174] = 8'd132;
   assign soundFileAmplitudes [6175] = 8'd120;
   assign soundFileAmplitudes [6176] = 8'd102;
   assign soundFileAmplitudes [6177] = 8'd96;
   assign soundFileAmplitudes [6178] = 8'd101;
   assign soundFileAmplitudes [6179] = 8'd117;
   assign soundFileAmplitudes [6180] = 8'd120;
   assign soundFileAmplitudes [6181] = 8'd116;
   assign soundFileAmplitudes [6182] = 8'd114;
   assign soundFileAmplitudes [6183] = 8'd123;
   assign soundFileAmplitudes [6184] = 8'd126;
   assign soundFileAmplitudes [6185] = 8'd134;
   assign soundFileAmplitudes [6186] = 8'd144;
   assign soundFileAmplitudes [6187] = 8'd140;
   assign soundFileAmplitudes [6188] = 8'd141;
   assign soundFileAmplitudes [6189] = 8'd131;
   assign soundFileAmplitudes [6190] = 8'd125;
   assign soundFileAmplitudes [6191] = 8'd123;
   assign soundFileAmplitudes [6192] = 8'd113;
   assign soundFileAmplitudes [6193] = 8'd111;
   assign soundFileAmplitudes [6194] = 8'd110;
   assign soundFileAmplitudes [6195] = 8'd116;
   assign soundFileAmplitudes [6196] = 8'd116;
   assign soundFileAmplitudes [6197] = 8'd121;
   assign soundFileAmplitudes [6198] = 8'd118;
   assign soundFileAmplitudes [6199] = 8'd118;
   assign soundFileAmplitudes [6200] = 8'd133;
   assign soundFileAmplitudes [6201] = 8'd138;
   assign soundFileAmplitudes [6202] = 8'd145;
   assign soundFileAmplitudes [6203] = 8'd149;
   assign soundFileAmplitudes [6204] = 8'd142;
   assign soundFileAmplitudes [6205] = 8'd132;
   assign soundFileAmplitudes [6206] = 8'd139;
   assign soundFileAmplitudes [6207] = 8'd134;
   assign soundFileAmplitudes [6208] = 8'd124;
   assign soundFileAmplitudes [6209] = 8'd120;
   assign soundFileAmplitudes [6210] = 8'd125;
   assign soundFileAmplitudes [6211] = 8'd120;
   assign soundFileAmplitudes [6212] = 8'd96;
   assign soundFileAmplitudes [6213] = 8'd92;
   assign soundFileAmplitudes [6214] = 8'd92;
   assign soundFileAmplitudes [6215] = 8'd114;
   assign soundFileAmplitudes [6216] = 8'd136;
   assign soundFileAmplitudes [6217] = 8'd133;
   assign soundFileAmplitudes [6218] = 8'd126;
   assign soundFileAmplitudes [6219] = 8'd125;
   assign soundFileAmplitudes [6220] = 8'd133;
   assign soundFileAmplitudes [6221] = 8'd147;
   assign soundFileAmplitudes [6222] = 8'd158;
   assign soundFileAmplitudes [6223] = 8'd154;
   assign soundFileAmplitudes [6224] = 8'd137;
   assign soundFileAmplitudes [6225] = 8'd116;
   assign soundFileAmplitudes [6226] = 8'd110;
   assign soundFileAmplitudes [6227] = 8'd105;
   assign soundFileAmplitudes [6228] = 8'd109;
   assign soundFileAmplitudes [6229] = 8'd120;
   assign soundFileAmplitudes [6230] = 8'd124;
   assign soundFileAmplitudes [6231] = 8'd123;
   assign soundFileAmplitudes [6232] = 8'd118;
   assign soundFileAmplitudes [6233] = 8'd112;
   assign soundFileAmplitudes [6234] = 8'd114;
   assign soundFileAmplitudes [6235] = 8'd124;
   assign soundFileAmplitudes [6236] = 8'd135;
   assign soundFileAmplitudes [6237] = 8'd151;
   assign soundFileAmplitudes [6238] = 8'd154;
   assign soundFileAmplitudes [6239] = 8'd150;
   assign soundFileAmplitudes [6240] = 8'd138;
   assign soundFileAmplitudes [6241] = 8'd127;
   assign soundFileAmplitudes [6242] = 8'd130;
   assign soundFileAmplitudes [6243] = 8'd130;
   assign soundFileAmplitudes [6244] = 8'd126;
   assign soundFileAmplitudes [6245] = 8'd120;
   assign soundFileAmplitudes [6246] = 8'd111;
   assign soundFileAmplitudes [6247] = 8'd97;
   assign soundFileAmplitudes [6248] = 8'd89;
   assign soundFileAmplitudes [6249] = 8'd93;
   assign soundFileAmplitudes [6250] = 8'd107;
   assign soundFileAmplitudes [6251] = 8'd126;
   assign soundFileAmplitudes [6252] = 8'd134;
   assign soundFileAmplitudes [6253] = 8'd132;
   assign soundFileAmplitudes [6254] = 8'd131;
   assign soundFileAmplitudes [6255] = 8'd136;
   assign soundFileAmplitudes [6256] = 8'd152;
   assign soundFileAmplitudes [6257] = 8'd159;
   assign soundFileAmplitudes [6258] = 8'd148;
   assign soundFileAmplitudes [6259] = 8'd145;
   assign soundFileAmplitudes [6260] = 8'd136;
   assign soundFileAmplitudes [6261] = 8'd124;
   assign soundFileAmplitudes [6262] = 8'd117;
   assign soundFileAmplitudes [6263] = 8'd109;
   assign soundFileAmplitudes [6264] = 8'd104;
   assign soundFileAmplitudes [6265] = 8'd103;
   assign soundFileAmplitudes [6266] = 8'd107;
   assign soundFileAmplitudes [6267] = 8'd101;
   assign soundFileAmplitudes [6268] = 8'd100;
   assign soundFileAmplitudes [6269] = 8'd112;
   assign soundFileAmplitudes [6270] = 8'd121;
   assign soundFileAmplitudes [6271] = 8'd136;
   assign soundFileAmplitudes [6272] = 8'd142;
   assign soundFileAmplitudes [6273] = 8'd147;
   assign soundFileAmplitudes [6274] = 8'd143;
   assign soundFileAmplitudes [6275] = 8'd132;
   assign soundFileAmplitudes [6276] = 8'd136;
   assign soundFileAmplitudes [6277] = 8'd138;
   assign soundFileAmplitudes [6278] = 8'd145;
   assign soundFileAmplitudes [6279] = 8'd151;
   assign soundFileAmplitudes [6280] = 8'd145;
   assign soundFileAmplitudes [6281] = 8'd127;
   assign soundFileAmplitudes [6282] = 8'd115;
   assign soundFileAmplitudes [6283] = 8'd102;
   assign soundFileAmplitudes [6284] = 8'd108;
   assign soundFileAmplitudes [6285] = 8'd127;
   assign soundFileAmplitudes [6286] = 8'd141;
   assign soundFileAmplitudes [6287] = 8'd138;
   assign soundFileAmplitudes [6288] = 8'd126;
   assign soundFileAmplitudes [6289] = 8'd124;
   assign soundFileAmplitudes [6290] = 8'd129;
   assign soundFileAmplitudes [6291] = 8'd146;
   assign soundFileAmplitudes [6292] = 8'd157;
   assign soundFileAmplitudes [6293] = 8'd148;
   assign soundFileAmplitudes [6294] = 8'd137;
   assign soundFileAmplitudes [6295] = 8'd135;
   assign soundFileAmplitudes [6296] = 8'd132;
   assign soundFileAmplitudes [6297] = 8'd123;
   assign soundFileAmplitudes [6298] = 8'd108;
   assign soundFileAmplitudes [6299] = 8'd105;
   assign soundFileAmplitudes [6300] = 8'd113;
   assign soundFileAmplitudes [6301] = 8'd127;
   assign soundFileAmplitudes [6302] = 8'd122;
   assign soundFileAmplitudes [6303] = 8'd111;
   assign soundFileAmplitudes [6304] = 8'd109;
   assign soundFileAmplitudes [6305] = 8'd113;
   assign soundFileAmplitudes [6306] = 8'd125;
   assign soundFileAmplitudes [6307] = 8'd128;
   assign soundFileAmplitudes [6308] = 8'd138;
   assign soundFileAmplitudes [6309] = 8'd131;
   assign soundFileAmplitudes [6310] = 8'd125;
   assign soundFileAmplitudes [6311] = 8'd124;
   assign soundFileAmplitudes [6312] = 8'd122;
   assign soundFileAmplitudes [6313] = 8'd128;
   assign soundFileAmplitudes [6314] = 8'd130;
   assign soundFileAmplitudes [6315] = 8'd125;
   assign soundFileAmplitudes [6316] = 8'd122;
   assign soundFileAmplitudes [6317] = 8'd112;
   assign soundFileAmplitudes [6318] = 8'd93;
   assign soundFileAmplitudes [6319] = 8'd87;
   assign soundFileAmplitudes [6320] = 8'd113;
   assign soundFileAmplitudes [6321] = 8'd142;
   assign soundFileAmplitudes [6322] = 8'd145;
   assign soundFileAmplitudes [6323] = 8'd130;
   assign soundFileAmplitudes [6324] = 8'd117;
   assign soundFileAmplitudes [6325] = 8'd120;
   assign soundFileAmplitudes [6326] = 8'd145;
   assign soundFileAmplitudes [6327] = 8'd152;
   assign soundFileAmplitudes [6328] = 8'd144;
   assign soundFileAmplitudes [6329] = 8'd147;
   assign soundFileAmplitudes [6330] = 8'd123;
   assign soundFileAmplitudes [6331] = 8'd119;
   assign soundFileAmplitudes [6332] = 8'd118;
   assign soundFileAmplitudes [6333] = 8'd118;
   assign soundFileAmplitudes [6334] = 8'd119;
   assign soundFileAmplitudes [6335] = 8'd110;
   assign soundFileAmplitudes [6336] = 8'd115;
   assign soundFileAmplitudes [6337] = 8'd111;
   assign soundFileAmplitudes [6338] = 8'd118;
   assign soundFileAmplitudes [6339] = 8'd122;
   assign soundFileAmplitudes [6340] = 8'd133;
   assign soundFileAmplitudes [6341] = 8'd142;
   assign soundFileAmplitudes [6342] = 8'd152;
   assign soundFileAmplitudes [6343] = 8'd155;
   assign soundFileAmplitudes [6344] = 8'd149;
   assign soundFileAmplitudes [6345] = 8'd146;
   assign soundFileAmplitudes [6346] = 8'd130;
   assign soundFileAmplitudes [6347] = 8'd128;
   assign soundFileAmplitudes [6348] = 8'd131;
   assign soundFileAmplitudes [6349] = 8'd127;
   assign soundFileAmplitudes [6350] = 8'd125;
   assign soundFileAmplitudes [6351] = 8'd129;
   assign soundFileAmplitudes [6352] = 8'd111;
   assign soundFileAmplitudes [6353] = 8'd88;
   assign soundFileAmplitudes [6354] = 8'd90;
   assign soundFileAmplitudes [6355] = 8'd104;
   assign soundFileAmplitudes [6356] = 8'd122;
   assign soundFileAmplitudes [6357] = 8'd124;
   assign soundFileAmplitudes [6358] = 8'd115;
   assign soundFileAmplitudes [6359] = 8'd109;
   assign soundFileAmplitudes [6360] = 8'd120;
   assign soundFileAmplitudes [6361] = 8'd136;
   assign soundFileAmplitudes [6362] = 8'd139;
   assign soundFileAmplitudes [6363] = 8'd139;
   assign soundFileAmplitudes [6364] = 8'd139;
   assign soundFileAmplitudes [6365] = 8'd124;
   assign soundFileAmplitudes [6366] = 8'd113;
   assign soundFileAmplitudes [6367] = 8'd110;
   assign soundFileAmplitudes [6368] = 8'd107;
   assign soundFileAmplitudes [6369] = 8'd122;
   assign soundFileAmplitudes [6370] = 8'd127;
   assign soundFileAmplitudes [6371] = 8'd129;
   assign soundFileAmplitudes [6372] = 8'd129;
   assign soundFileAmplitudes [6373] = 8'd128;
   assign soundFileAmplitudes [6374] = 8'd126;
   assign soundFileAmplitudes [6375] = 8'd125;
   assign soundFileAmplitudes [6376] = 8'd139;
   assign soundFileAmplitudes [6377] = 8'd150;
   assign soundFileAmplitudes [6378] = 8'd160;
   assign soundFileAmplitudes [6379] = 8'd158;
   assign soundFileAmplitudes [6380] = 8'd147;
   assign soundFileAmplitudes [6381] = 8'd139;
   assign soundFileAmplitudes [6382] = 8'd136;
   assign soundFileAmplitudes [6383] = 8'd135;
   assign soundFileAmplitudes [6384] = 8'd134;
   assign soundFileAmplitudes [6385] = 8'd129;
   assign soundFileAmplitudes [6386] = 8'd117;
   assign soundFileAmplitudes [6387] = 8'd107;
   assign soundFileAmplitudes [6388] = 8'd89;
   assign soundFileAmplitudes [6389] = 8'd78;
   assign soundFileAmplitudes [6390] = 8'd90;
   assign soundFileAmplitudes [6391] = 8'd108;
   assign soundFileAmplitudes [6392] = 8'd115;
   assign soundFileAmplitudes [6393] = 8'd116;
   assign soundFileAmplitudes [6394] = 8'd116;
   assign soundFileAmplitudes [6395] = 8'd124;
   assign soundFileAmplitudes [6396] = 8'd145;
   assign soundFileAmplitudes [6397] = 8'd147;
   assign soundFileAmplitudes [6398] = 8'd145;
   assign soundFileAmplitudes [6399] = 8'd145;
   assign soundFileAmplitudes [6400] = 8'd132;
   assign soundFileAmplitudes [6401] = 8'd133;
   assign soundFileAmplitudes [6402] = 8'd130;
   assign soundFileAmplitudes [6403] = 8'd130;
   assign soundFileAmplitudes [6404] = 8'd129;
   assign soundFileAmplitudes [6405] = 8'd133;
   assign soundFileAmplitudes [6406] = 8'd132;
   assign soundFileAmplitudes [6407] = 8'd123;
   assign soundFileAmplitudes [6408] = 8'd120;
   assign soundFileAmplitudes [6409] = 8'd115;
   assign soundFileAmplitudes [6410] = 8'd116;
   assign soundFileAmplitudes [6411] = 8'd116;
   assign soundFileAmplitudes [6412] = 8'd123;
   assign soundFileAmplitudes [6413] = 8'd132;
   assign soundFileAmplitudes [6414] = 8'd140;
   assign soundFileAmplitudes [6415] = 8'd138;
   assign soundFileAmplitudes [6416] = 8'd132;
   assign soundFileAmplitudes [6417] = 8'd131;
   assign soundFileAmplitudes [6418] = 8'd132;
   assign soundFileAmplitudes [6419] = 8'd138;
   assign soundFileAmplitudes [6420] = 8'd133;
   assign soundFileAmplitudes [6421] = 8'd122;
   assign soundFileAmplitudes [6422] = 8'd114;
   assign soundFileAmplitudes [6423] = 8'd101;
   assign soundFileAmplitudes [6424] = 8'd97;
   assign soundFileAmplitudes [6425] = 8'd116;
   assign soundFileAmplitudes [6426] = 8'd128;
   assign soundFileAmplitudes [6427] = 8'd128;
   assign soundFileAmplitudes [6428] = 8'd120;
   assign soundFileAmplitudes [6429] = 8'd122;
   assign soundFileAmplitudes [6430] = 8'd129;
   assign soundFileAmplitudes [6431] = 8'd144;
   assign soundFileAmplitudes [6432] = 8'd153;
   assign soundFileAmplitudes [6433] = 8'd148;
   assign soundFileAmplitudes [6434] = 8'd149;
   assign soundFileAmplitudes [6435] = 8'd141;
   assign soundFileAmplitudes [6436] = 8'd140;
   assign soundFileAmplitudes [6437] = 8'd135;
   assign soundFileAmplitudes [6438] = 8'd123;
   assign soundFileAmplitudes [6439] = 8'd120;
   assign soundFileAmplitudes [6440] = 8'd123;
   assign soundFileAmplitudes [6441] = 8'd124;
   assign soundFileAmplitudes [6442] = 8'd120;
   assign soundFileAmplitudes [6443] = 8'd113;
   assign soundFileAmplitudes [6444] = 8'd112;
   assign soundFileAmplitudes [6445] = 8'd113;
   assign soundFileAmplitudes [6446] = 8'd118;
   assign soundFileAmplitudes [6447] = 8'd119;
   assign soundFileAmplitudes [6448] = 8'd123;
   assign soundFileAmplitudes [6449] = 8'd127;
   assign soundFileAmplitudes [6450] = 8'd132;
   assign soundFileAmplitudes [6451] = 8'd134;
   assign soundFileAmplitudes [6452] = 8'd127;
   assign soundFileAmplitudes [6453] = 8'd133;
   assign soundFileAmplitudes [6454] = 8'd133;
   assign soundFileAmplitudes [6455] = 8'd123;
   assign soundFileAmplitudes [6456] = 8'd118;
   assign soundFileAmplitudes [6457] = 8'd105;
   assign soundFileAmplitudes [6458] = 8'd94;
   assign soundFileAmplitudes [6459] = 8'd90;
   assign soundFileAmplitudes [6460] = 8'd98;
   assign soundFileAmplitudes [6461] = 8'd115;
   assign soundFileAmplitudes [6462] = 8'd124;
   assign soundFileAmplitudes [6463] = 8'd131;
   assign soundFileAmplitudes [6464] = 8'd130;
   assign soundFileAmplitudes [6465] = 8'd123;
   assign soundFileAmplitudes [6466] = 8'd142;
   assign soundFileAmplitudes [6467] = 8'd171;
   assign soundFileAmplitudes [6468] = 8'd162;
   assign soundFileAmplitudes [6469] = 8'd160;
   assign soundFileAmplitudes [6470] = 8'd158;
   assign soundFileAmplitudes [6471] = 8'd155;
   assign soundFileAmplitudes [6472] = 8'd153;
   assign soundFileAmplitudes [6473] = 8'd144;
   assign soundFileAmplitudes [6474] = 8'd135;
   assign soundFileAmplitudes [6475] = 8'd126;
   assign soundFileAmplitudes [6476] = 8'd126;
   assign soundFileAmplitudes [6477] = 8'd114;
   assign soundFileAmplitudes [6478] = 8'd108;
   assign soundFileAmplitudes [6479] = 8'd101;
   assign soundFileAmplitudes [6480] = 8'd97;
   assign soundFileAmplitudes [6481] = 8'd107;
   assign soundFileAmplitudes [6482] = 8'd114;
   assign soundFileAmplitudes [6483] = 8'd117;
   assign soundFileAmplitudes [6484] = 8'd118;
   assign soundFileAmplitudes [6485] = 8'd116;
   assign soundFileAmplitudes [6486] = 8'd120;
   assign soundFileAmplitudes [6487] = 8'd119;
   assign soundFileAmplitudes [6488] = 8'd125;
   assign soundFileAmplitudes [6489] = 8'd127;
   assign soundFileAmplitudes [6490] = 8'd122;
   assign soundFileAmplitudes [6491] = 8'd107;
   assign soundFileAmplitudes [6492] = 8'd101;
   assign soundFileAmplitudes [6493] = 8'd93;
   assign soundFileAmplitudes [6494] = 8'd84;
   assign soundFileAmplitudes [6495] = 8'd99;
   assign soundFileAmplitudes [6496] = 8'd116;
   assign soundFileAmplitudes [6497] = 8'd125;
   assign soundFileAmplitudes [6498] = 8'd131;
   assign soundFileAmplitudes [6499] = 8'd134;
   assign soundFileAmplitudes [6500] = 8'd139;
   assign soundFileAmplitudes [6501] = 8'd143;
   assign soundFileAmplitudes [6502] = 8'd154;
   assign soundFileAmplitudes [6503] = 8'd168;
   assign soundFileAmplitudes [6504] = 8'd166;
   assign soundFileAmplitudes [6505] = 8'd172;
   assign soundFileAmplitudes [6506] = 8'd166;
   assign soundFileAmplitudes [6507] = 8'd153;
   assign soundFileAmplitudes [6508] = 8'd137;
   assign soundFileAmplitudes [6509] = 8'd128;
   assign soundFileAmplitudes [6510] = 8'd127;
   assign soundFileAmplitudes [6511] = 8'd127;
   assign soundFileAmplitudes [6512] = 8'd130;
   assign soundFileAmplitudes [6513] = 8'd119;
   assign soundFileAmplitudes [6514] = 8'd110;
   assign soundFileAmplitudes [6515] = 8'd107;
   assign soundFileAmplitudes [6516] = 8'd103;
   assign soundFileAmplitudes [6517] = 8'd105;
   assign soundFileAmplitudes [6518] = 8'd113;
   assign soundFileAmplitudes [6519] = 8'd119;
   assign soundFileAmplitudes [6520] = 8'd124;
   assign soundFileAmplitudes [6521] = 8'd116;
   assign soundFileAmplitudes [6522] = 8'd119;
   assign soundFileAmplitudes [6523] = 8'd116;
   assign soundFileAmplitudes [6524] = 8'd117;
   assign soundFileAmplitudes [6525] = 8'd124;
   assign soundFileAmplitudes [6526] = 8'd120;
   assign soundFileAmplitudes [6527] = 8'd120;
   assign soundFileAmplitudes [6528] = 8'd119;
   assign soundFileAmplitudes [6529] = 8'd116;
   assign soundFileAmplitudes [6530] = 8'd105;
   assign soundFileAmplitudes [6531] = 8'd102;
   assign soundFileAmplitudes [6532] = 8'd116;
   assign soundFileAmplitudes [6533] = 8'd132;
   assign soundFileAmplitudes [6534] = 8'd141;
   assign soundFileAmplitudes [6535] = 8'd145;
   assign soundFileAmplitudes [6536] = 8'd136;
   assign soundFileAmplitudes [6537] = 8'd131;
   assign soundFileAmplitudes [6538] = 8'd141;
   assign soundFileAmplitudes [6539] = 8'd155;
   assign soundFileAmplitudes [6540] = 8'd158;
   assign soundFileAmplitudes [6541] = 8'd162;
   assign soundFileAmplitudes [6542] = 8'd153;
   assign soundFileAmplitudes [6543] = 8'd136;
   assign soundFileAmplitudes [6544] = 8'd116;
   assign soundFileAmplitudes [6545] = 8'd112;
   assign soundFileAmplitudes [6546] = 8'd121;
   assign soundFileAmplitudes [6547] = 8'd132;
   assign soundFileAmplitudes [6548] = 8'd140;
   assign soundFileAmplitudes [6549] = 8'd135;
   assign soundFileAmplitudes [6550] = 8'd121;
   assign soundFileAmplitudes [6551] = 8'd104;
   assign soundFileAmplitudes [6552] = 8'd107;
   assign soundFileAmplitudes [6553] = 8'd108;
   assign soundFileAmplitudes [6554] = 8'd117;
   assign soundFileAmplitudes [6555] = 8'd121;
   assign soundFileAmplitudes [6556] = 8'd125;
   assign soundFileAmplitudes [6557] = 8'd130;
   assign soundFileAmplitudes [6558] = 8'd123;
   assign soundFileAmplitudes [6559] = 8'd119;
   assign soundFileAmplitudes [6560] = 8'd123;
   assign soundFileAmplitudes [6561] = 8'd124;
   assign soundFileAmplitudes [6562] = 8'd116;
   assign soundFileAmplitudes [6563] = 8'd117;
   assign soundFileAmplitudes [6564] = 8'd121;
   assign soundFileAmplitudes [6565] = 8'd106;
   assign soundFileAmplitudes [6566] = 8'd99;
   assign soundFileAmplitudes [6567] = 8'd112;
   assign soundFileAmplitudes [6568] = 8'd129;
   assign soundFileAmplitudes [6569] = 8'd146;
   assign soundFileAmplitudes [6570] = 8'd151;
   assign soundFileAmplitudes [6571] = 8'd150;
   assign soundFileAmplitudes [6572] = 8'd139;
   assign soundFileAmplitudes [6573] = 8'd139;
   assign soundFileAmplitudes [6574] = 8'd153;
   assign soundFileAmplitudes [6575] = 8'd167;
   assign soundFileAmplitudes [6576] = 8'd158;
   assign soundFileAmplitudes [6577] = 8'd148;
   assign soundFileAmplitudes [6578] = 8'd143;
   assign soundFileAmplitudes [6579] = 8'd135;
   assign soundFileAmplitudes [6580] = 8'd119;
   assign soundFileAmplitudes [6581] = 8'd108;
   assign soundFileAmplitudes [6582] = 8'd111;
   assign soundFileAmplitudes [6583] = 8'd110;
   assign soundFileAmplitudes [6584] = 8'd106;
   assign soundFileAmplitudes [6585] = 8'd101;
   assign soundFileAmplitudes [6586] = 8'd98;
   assign soundFileAmplitudes [6587] = 8'd91;
   assign soundFileAmplitudes [6588] = 8'd98;
   assign soundFileAmplitudes [6589] = 8'd105;
   assign soundFileAmplitudes [6590] = 8'd117;
   assign soundFileAmplitudes [6591] = 8'd127;
   assign soundFileAmplitudes [6592] = 8'd141;
   assign soundFileAmplitudes [6593] = 8'd148;
   assign soundFileAmplitudes [6594] = 8'd148;
   assign soundFileAmplitudes [6595] = 8'd144;
   assign soundFileAmplitudes [6596] = 8'd142;
   assign soundFileAmplitudes [6597] = 8'd144;
   assign soundFileAmplitudes [6598] = 8'd139;
   assign soundFileAmplitudes [6599] = 8'd133;
   assign soundFileAmplitudes [6600] = 8'd122;
   assign soundFileAmplitudes [6601] = 8'd112;
   assign soundFileAmplitudes [6602] = 8'd101;
   assign soundFileAmplitudes [6603] = 8'd99;
   assign soundFileAmplitudes [6604] = 8'd107;
   assign soundFileAmplitudes [6605] = 8'd125;
   assign soundFileAmplitudes [6606] = 8'd132;
   assign soundFileAmplitudes [6607] = 8'd135;
   assign soundFileAmplitudes [6608] = 8'd138;
   assign soundFileAmplitudes [6609] = 8'd133;
   assign soundFileAmplitudes [6610] = 8'd130;
   assign soundFileAmplitudes [6611] = 8'd134;
   assign soundFileAmplitudes [6612] = 8'd141;
   assign soundFileAmplitudes [6613] = 8'd143;
   assign soundFileAmplitudes [6614] = 8'd140;
   assign soundFileAmplitudes [6615] = 8'd140;
   assign soundFileAmplitudes [6616] = 8'd131;
   assign soundFileAmplitudes [6617] = 8'd106;
   assign soundFileAmplitudes [6618] = 8'd102;
   assign soundFileAmplitudes [6619] = 8'd107;
   assign soundFileAmplitudes [6620] = 8'd113;
   assign soundFileAmplitudes [6621] = 8'd114;
   assign soundFileAmplitudes [6622] = 8'd111;
   assign soundFileAmplitudes [6623] = 8'd110;
   assign soundFileAmplitudes [6624] = 8'd118;
   assign soundFileAmplitudes [6625] = 8'd117;
   assign soundFileAmplitudes [6626] = 8'd122;
   assign soundFileAmplitudes [6627] = 8'd139;
   assign soundFileAmplitudes [6628] = 8'd143;
   assign soundFileAmplitudes [6629] = 8'd146;
   assign soundFileAmplitudes [6630] = 8'd140;
   assign soundFileAmplitudes [6631] = 8'd143;
   assign soundFileAmplitudes [6632] = 8'd137;
   assign soundFileAmplitudes [6633] = 8'd131;
   assign soundFileAmplitudes [6634] = 8'd130;
   assign soundFileAmplitudes [6635] = 8'd122;
   assign soundFileAmplitudes [6636] = 8'd121;
   assign soundFileAmplitudes [6637] = 8'd116;
   assign soundFileAmplitudes [6638] = 8'd103;
   assign soundFileAmplitudes [6639] = 8'd98;
   assign soundFileAmplitudes [6640] = 8'd100;
   assign soundFileAmplitudes [6641] = 8'd111;
   assign soundFileAmplitudes [6642] = 8'd124;
   assign soundFileAmplitudes [6643] = 8'd127;
   assign soundFileAmplitudes [6644] = 8'd125;
   assign soundFileAmplitudes [6645] = 8'd125;
   assign soundFileAmplitudes [6646] = 8'd126;
   assign soundFileAmplitudes [6647] = 8'd127;
   assign soundFileAmplitudes [6648] = 8'd141;
   assign soundFileAmplitudes [6649] = 8'd155;
   assign soundFileAmplitudes [6650] = 8'd152;
   assign soundFileAmplitudes [6651] = 8'd144;
   assign soundFileAmplitudes [6652] = 8'd141;
   assign soundFileAmplitudes [6653] = 8'd141;
   assign soundFileAmplitudes [6654] = 8'd130;
   assign soundFileAmplitudes [6655] = 8'd118;
   assign soundFileAmplitudes [6656] = 8'd117;
   assign soundFileAmplitudes [6657] = 8'd121;
   assign soundFileAmplitudes [6658] = 8'd124;
   assign soundFileAmplitudes [6659] = 8'd117;
   assign soundFileAmplitudes [6660] = 8'd113;
   assign soundFileAmplitudes [6661] = 8'd114;
   assign soundFileAmplitudes [6662] = 8'd119;
   assign soundFileAmplitudes [6663] = 8'd125;
   assign soundFileAmplitudes [6664] = 8'd132;
   assign soundFileAmplitudes [6665] = 8'd132;
   assign soundFileAmplitudes [6666] = 8'd140;
   assign soundFileAmplitudes [6667] = 8'd136;
   assign soundFileAmplitudes [6668] = 8'd131;
   assign soundFileAmplitudes [6669] = 8'd130;
   assign soundFileAmplitudes [6670] = 8'd124;
   assign soundFileAmplitudes [6671] = 8'd127;
   assign soundFileAmplitudes [6672] = 8'd121;
   assign soundFileAmplitudes [6673] = 8'd113;
   assign soundFileAmplitudes [6674] = 8'd105;
   assign soundFileAmplitudes [6675] = 8'd96;
   assign soundFileAmplitudes [6676] = 8'd88;
   assign soundFileAmplitudes [6677] = 8'd89;
   assign soundFileAmplitudes [6678] = 8'd101;
   assign soundFileAmplitudes [6679] = 8'd116;
   assign soundFileAmplitudes [6680] = 8'd132;
   assign soundFileAmplitudes [6681] = 8'd145;
   assign soundFileAmplitudes [6682] = 8'd154;
   assign soundFileAmplitudes [6683] = 8'd153;
   assign soundFileAmplitudes [6684] = 8'd150;
   assign soundFileAmplitudes [6685] = 8'd150;
   assign soundFileAmplitudes [6686] = 8'd165;
   assign soundFileAmplitudes [6687] = 8'd159;
   assign soundFileAmplitudes [6688] = 8'd153;
   assign soundFileAmplitudes [6689] = 8'd151;
   assign soundFileAmplitudes [6690] = 8'd138;
   assign soundFileAmplitudes [6691] = 8'd137;
   assign soundFileAmplitudes [6692] = 8'd115;
   assign soundFileAmplitudes [6693] = 8'd110;
   assign soundFileAmplitudes [6694] = 8'd113;
   assign soundFileAmplitudes [6695] = 8'd123;
   assign soundFileAmplitudes [6696] = 8'd131;
   assign soundFileAmplitudes [6697] = 8'd122;
   assign soundFileAmplitudes [6698] = 8'd113;
   assign soundFileAmplitudes [6699] = 8'd101;
   assign soundFileAmplitudes [6700] = 8'd107;
   assign soundFileAmplitudes [6701] = 8'd119;
   assign soundFileAmplitudes [6702] = 8'd136;
   assign soundFileAmplitudes [6703] = 8'd144;
   assign soundFileAmplitudes [6704] = 8'd146;
   assign soundFileAmplitudes [6705] = 8'd140;
   assign soundFileAmplitudes [6706] = 8'd128;
   assign soundFileAmplitudes [6707] = 8'd122;
   assign soundFileAmplitudes [6708] = 8'd118;
   assign soundFileAmplitudes [6709] = 8'd112;
   assign soundFileAmplitudes [6710] = 8'd113;
   assign soundFileAmplitudes [6711] = 8'd116;
   assign soundFileAmplitudes [6712] = 8'd112;
   assign soundFileAmplitudes [6713] = 8'd98;
   assign soundFileAmplitudes [6714] = 8'd85;
   assign soundFileAmplitudes [6715] = 8'd94;
   assign soundFileAmplitudes [6716] = 8'd103;
   assign soundFileAmplitudes [6717] = 8'd117;
   assign soundFileAmplitudes [6718] = 8'd132;
   assign soundFileAmplitudes [6719] = 8'd150;
   assign soundFileAmplitudes [6720] = 8'd153;
   assign soundFileAmplitudes [6721] = 8'd144;
   assign soundFileAmplitudes [6722] = 8'd144;
   assign soundFileAmplitudes [6723] = 8'd153;
   assign soundFileAmplitudes [6724] = 8'd156;
   assign soundFileAmplitudes [6725] = 8'd156;
   assign soundFileAmplitudes [6726] = 8'd157;
   assign soundFileAmplitudes [6727] = 8'd149;
   assign soundFileAmplitudes [6728] = 8'd148;
   assign soundFileAmplitudes [6729] = 8'd127;
   assign soundFileAmplitudes [6730] = 8'd103;
   assign soundFileAmplitudes [6731] = 8'd107;
   assign soundFileAmplitudes [6732] = 8'd113;
   assign soundFileAmplitudes [6733] = 8'd116;
   assign soundFileAmplitudes [6734] = 8'd116;
   assign soundFileAmplitudes [6735] = 8'd112;
   assign soundFileAmplitudes [6736] = 8'd111;
   assign soundFileAmplitudes [6737] = 8'd108;
   assign soundFileAmplitudes [6738] = 8'd109;
   assign soundFileAmplitudes [6739] = 8'd132;
   assign soundFileAmplitudes [6740] = 8'd142;
   assign soundFileAmplitudes [6741] = 8'd143;
   assign soundFileAmplitudes [6742] = 8'd141;
   assign soundFileAmplitudes [6743] = 8'd132;
   assign soundFileAmplitudes [6744] = 8'd127;
   assign soundFileAmplitudes [6745] = 8'd121;
   assign soundFileAmplitudes [6746] = 8'd118;
   assign soundFileAmplitudes [6747] = 8'd120;
   assign soundFileAmplitudes [6748] = 8'd120;
   assign soundFileAmplitudes [6749] = 8'd118;
   assign soundFileAmplitudes [6750] = 8'd112;
   assign soundFileAmplitudes [6751] = 8'd104;
   assign soundFileAmplitudes [6752] = 8'd100;
   assign soundFileAmplitudes [6753] = 8'd101;
   assign soundFileAmplitudes [6754] = 8'd118;
   assign soundFileAmplitudes [6755] = 8'd129;
   assign soundFileAmplitudes [6756] = 8'd138;
   assign soundFileAmplitudes [6757] = 8'd139;
   assign soundFileAmplitudes [6758] = 8'd132;
   assign soundFileAmplitudes [6759] = 8'd131;
   assign soundFileAmplitudes [6760] = 8'd136;
   assign soundFileAmplitudes [6761] = 8'd147;
   assign soundFileAmplitudes [6762] = 8'd151;
   assign soundFileAmplitudes [6763] = 8'd146;
   assign soundFileAmplitudes [6764] = 8'd145;
   assign soundFileAmplitudes [6765] = 8'd145;
   assign soundFileAmplitudes [6766] = 8'd144;
   assign soundFileAmplitudes [6767] = 8'd122;
   assign soundFileAmplitudes [6768] = 8'd106;
   assign soundFileAmplitudes [6769] = 8'd107;
   assign soundFileAmplitudes [6770] = 8'd105;
   assign soundFileAmplitudes [6771] = 8'd117;
   assign soundFileAmplitudes [6772] = 8'd116;
   assign soundFileAmplitudes [6773] = 8'd111;
   assign soundFileAmplitudes [6774] = 8'd107;
   assign soundFileAmplitudes [6775] = 8'd105;
   assign soundFileAmplitudes [6776] = 8'd110;
   assign soundFileAmplitudes [6777] = 8'd128;
   assign soundFileAmplitudes [6778] = 8'd142;
   assign soundFileAmplitudes [6779] = 8'd149;
   assign soundFileAmplitudes [6780] = 8'd156;
   assign soundFileAmplitudes [6781] = 8'd153;
   assign soundFileAmplitudes [6782] = 8'd145;
   assign soundFileAmplitudes [6783] = 8'd132;
   assign soundFileAmplitudes [6784] = 8'd135;
   assign soundFileAmplitudes [6785] = 8'd131;
   assign soundFileAmplitudes [6786] = 8'd126;
   assign soundFileAmplitudes [6787] = 8'd126;
   assign soundFileAmplitudes [6788] = 8'd118;
   assign soundFileAmplitudes [6789] = 8'd102;
   assign soundFileAmplitudes [6790] = 8'd82;
   assign soundFileAmplitudes [6791] = 8'd78;
   assign soundFileAmplitudes [6792] = 8'd86;
   assign soundFileAmplitudes [6793] = 8'd102;
   assign soundFileAmplitudes [6794] = 8'd122;
   assign soundFileAmplitudes [6795] = 8'd137;
   assign soundFileAmplitudes [6796] = 8'd135;
   assign soundFileAmplitudes [6797] = 8'd128;
   assign soundFileAmplitudes [6798] = 8'd124;
   assign soundFileAmplitudes [6799] = 8'd137;
   assign soundFileAmplitudes [6800] = 8'd155;
   assign soundFileAmplitudes [6801] = 8'd155;
   assign soundFileAmplitudes [6802] = 8'd159;
   assign soundFileAmplitudes [6803] = 8'd159;
   assign soundFileAmplitudes [6804] = 8'd164;
   assign soundFileAmplitudes [6805] = 8'd140;
   assign soundFileAmplitudes [6806] = 8'd112;
   assign soundFileAmplitudes [6807] = 8'd108;
   assign soundFileAmplitudes [6808] = 8'd113;
   assign soundFileAmplitudes [6809] = 8'd127;
   assign soundFileAmplitudes [6810] = 8'd122;
   assign soundFileAmplitudes [6811] = 8'd113;
   assign soundFileAmplitudes [6812] = 8'd100;
   assign soundFileAmplitudes [6813] = 8'd93;
   assign soundFileAmplitudes [6814] = 8'd100;
   assign soundFileAmplitudes [6815] = 8'd130;
   assign soundFileAmplitudes [6816] = 8'd150;
   assign soundFileAmplitudes [6817] = 8'd158;
   assign soundFileAmplitudes [6818] = 8'd162;
   assign soundFileAmplitudes [6819] = 8'd154;
   assign soundFileAmplitudes [6820] = 8'd150;
   assign soundFileAmplitudes [6821] = 8'd141;
   assign soundFileAmplitudes [6822] = 8'd136;
   assign soundFileAmplitudes [6823] = 8'd136;
   assign soundFileAmplitudes [6824] = 8'd129;
   assign soundFileAmplitudes [6825] = 8'd121;
   assign soundFileAmplitudes [6826] = 8'd116;
   assign soundFileAmplitudes [6827] = 8'd97;
   assign soundFileAmplitudes [6828] = 8'd79;
   assign soundFileAmplitudes [6829] = 8'd78;
   assign soundFileAmplitudes [6830] = 8'd93;
   assign soundFileAmplitudes [6831] = 8'd119;
   assign soundFileAmplitudes [6832] = 8'd134;
   assign soundFileAmplitudes [6833] = 8'd141;
   assign soundFileAmplitudes [6834] = 8'd136;
   assign soundFileAmplitudes [6835] = 8'd123;
   assign soundFileAmplitudes [6836] = 8'd136;
   assign soundFileAmplitudes [6837] = 8'd146;
   assign soundFileAmplitudes [6838] = 8'd144;
   assign soundFileAmplitudes [6839] = 8'd144;
   assign soundFileAmplitudes [6840] = 8'd144;
   assign soundFileAmplitudes [6841] = 8'd147;
   assign soundFileAmplitudes [6842] = 8'd119;
   assign soundFileAmplitudes [6843] = 8'd98;
   assign soundFileAmplitudes [6844] = 8'd101;
   assign soundFileAmplitudes [6845] = 8'd109;
   assign soundFileAmplitudes [6846] = 8'd118;
   assign soundFileAmplitudes [6847] = 8'd115;
   assign soundFileAmplitudes [6848] = 8'd113;
   assign soundFileAmplitudes [6849] = 8'd110;
   assign soundFileAmplitudes [6850] = 8'd107;
   assign soundFileAmplitudes [6851] = 8'd107;
   assign soundFileAmplitudes [6852] = 8'd132;
   assign soundFileAmplitudes [6853] = 8'd156;
   assign soundFileAmplitudes [6854] = 8'd164;
   assign soundFileAmplitudes [6855] = 8'd170;
   assign soundFileAmplitudes [6856] = 8'd165;
   assign soundFileAmplitudes [6857] = 8'd156;
   assign soundFileAmplitudes [6858] = 8'd152;
   assign soundFileAmplitudes [6859] = 8'd145;
   assign soundFileAmplitudes [6860] = 8'd138;
   assign soundFileAmplitudes [6861] = 8'd131;
   assign soundFileAmplitudes [6862] = 8'd120;
   assign soundFileAmplitudes [6863] = 8'd110;
   assign soundFileAmplitudes [6864] = 8'd94;
   assign soundFileAmplitudes [6865] = 8'd89;
   assign soundFileAmplitudes [6866] = 8'd96;
   assign soundFileAmplitudes [6867] = 8'd108;
   assign soundFileAmplitudes [6868] = 8'd123;
   assign soundFileAmplitudes [6869] = 8'd125;
   assign soundFileAmplitudes [6870] = 8'd124;
   assign soundFileAmplitudes [6871] = 8'd119;
   assign soundFileAmplitudes [6872] = 8'd113;
   assign soundFileAmplitudes [6873] = 8'd127;
   assign soundFileAmplitudes [6874] = 8'd137;
   assign soundFileAmplitudes [6875] = 8'd135;
   assign soundFileAmplitudes [6876] = 8'd135;
   assign soundFileAmplitudes [6877] = 8'd138;
   assign soundFileAmplitudes [6878] = 8'd130;
   assign soundFileAmplitudes [6879] = 8'd101;
   assign soundFileAmplitudes [6880] = 8'd85;
   assign soundFileAmplitudes [6881] = 8'd90;
   assign soundFileAmplitudes [6882] = 8'd107;
   assign soundFileAmplitudes [6883] = 8'd125;
   assign soundFileAmplitudes [6884] = 8'd134;
   assign soundFileAmplitudes [6885] = 8'd128;
   assign soundFileAmplitudes [6886] = 8'd119;
   assign soundFileAmplitudes [6887] = 8'd117;
   assign soundFileAmplitudes [6888] = 8'd128;
   assign soundFileAmplitudes [6889] = 8'd153;
   assign soundFileAmplitudes [6890] = 8'd171;
   assign soundFileAmplitudes [6891] = 8'd182;
   assign soundFileAmplitudes [6892] = 8'd176;
   assign soundFileAmplitudes [6893] = 8'd168;
   assign soundFileAmplitudes [6894] = 8'd147;
   assign soundFileAmplitudes [6895] = 8'd129;
   assign soundFileAmplitudes [6896] = 8'd127;
   assign soundFileAmplitudes [6897] = 8'd121;
   assign soundFileAmplitudes [6898] = 8'd118;
   assign soundFileAmplitudes [6899] = 8'd116;
   assign soundFileAmplitudes [6900] = 8'd104;
   assign soundFileAmplitudes [6901] = 8'd89;
   assign soundFileAmplitudes [6902] = 8'd87;
   assign soundFileAmplitudes [6903] = 8'd92;
   assign soundFileAmplitudes [6904] = 8'd106;
   assign soundFileAmplitudes [6905] = 8'd121;
   assign soundFileAmplitudes [6906] = 8'd133;
   assign soundFileAmplitudes [6907] = 8'd133;
   assign soundFileAmplitudes [6908] = 8'd128;
   assign soundFileAmplitudes [6909] = 8'd128;
   assign soundFileAmplitudes [6910] = 8'd138;
   assign soundFileAmplitudes [6911] = 8'd141;
   assign soundFileAmplitudes [6912] = 8'd136;
   assign soundFileAmplitudes [6913] = 8'd138;
   assign soundFileAmplitudes [6914] = 8'd140;
   assign soundFileAmplitudes [6915] = 8'd132;
   assign soundFileAmplitudes [6916] = 8'd104;
   assign soundFileAmplitudes [6917] = 8'd89;
   assign soundFileAmplitudes [6918] = 8'd93;
   assign soundFileAmplitudes [6919] = 8'd105;
   assign soundFileAmplitudes [6920] = 8'd113;
   assign soundFileAmplitudes [6921] = 8'd109;
   assign soundFileAmplitudes [6922] = 8'd110;
   assign soundFileAmplitudes [6923] = 8'd105;
   assign soundFileAmplitudes [6924] = 8'd108;
   assign soundFileAmplitudes [6925] = 8'd131;
   assign soundFileAmplitudes [6926] = 8'd151;
   assign soundFileAmplitudes [6927] = 8'd162;
   assign soundFileAmplitudes [6928] = 8'd168;
   assign soundFileAmplitudes [6929] = 8'd165;
   assign soundFileAmplitudes [6930] = 8'd159;
   assign soundFileAmplitudes [6931] = 8'd150;
   assign soundFileAmplitudes [6932] = 8'd146;
   assign soundFileAmplitudes [6933] = 8'd137;
   assign soundFileAmplitudes [6934] = 8'd125;
   assign soundFileAmplitudes [6935] = 8'd126;
   assign soundFileAmplitudes [6936] = 8'd117;
   assign soundFileAmplitudes [6937] = 8'd109;
   assign soundFileAmplitudes [6938] = 8'd98;
   assign soundFileAmplitudes [6939] = 8'd93;
   assign soundFileAmplitudes [6940] = 8'd112;
   assign soundFileAmplitudes [6941] = 8'd128;
   assign soundFileAmplitudes [6942] = 8'd139;
   assign soundFileAmplitudes [6943] = 8'd142;
   assign soundFileAmplitudes [6944] = 8'd135;
   assign soundFileAmplitudes [6945] = 8'd125;
   assign soundFileAmplitudes [6946] = 8'd128;
   assign soundFileAmplitudes [6947] = 8'd147;
   assign soundFileAmplitudes [6948] = 8'd148;
   assign soundFileAmplitudes [6949] = 8'd145;
   assign soundFileAmplitudes [6950] = 8'd143;
   assign soundFileAmplitudes [6951] = 8'd130;
   assign soundFileAmplitudes [6952] = 8'd104;
   assign soundFileAmplitudes [6953] = 8'd76;
   assign soundFileAmplitudes [6954] = 8'd72;
   assign soundFileAmplitudes [6955] = 8'd90;
   assign soundFileAmplitudes [6956] = 8'd108;
   assign soundFileAmplitudes [6957] = 8'd112;
   assign soundFileAmplitudes [6958] = 8'd108;
   assign soundFileAmplitudes [6959] = 8'd107;
   assign soundFileAmplitudes [6960] = 8'd112;
   assign soundFileAmplitudes [6961] = 8'd128;
   assign soundFileAmplitudes [6962] = 8'd152;
   assign soundFileAmplitudes [6963] = 8'd172;
   assign soundFileAmplitudes [6964] = 8'd187;
   assign soundFileAmplitudes [6965] = 8'd188;
   assign soundFileAmplitudes [6966] = 8'd175;
   assign soundFileAmplitudes [6967] = 8'd159;
   assign soundFileAmplitudes [6968] = 8'd148;
   assign soundFileAmplitudes [6969] = 8'd145;
   assign soundFileAmplitudes [6970] = 8'd135;
   assign soundFileAmplitudes [6971] = 8'd125;
   assign soundFileAmplitudes [6972] = 8'd124;
   assign soundFileAmplitudes [6973] = 8'd118;
   assign soundFileAmplitudes [6974] = 8'd107;
   assign soundFileAmplitudes [6975] = 8'd89;
   assign soundFileAmplitudes [6976] = 8'd91;
   assign soundFileAmplitudes [6977] = 8'd109;
   assign soundFileAmplitudes [6978] = 8'd121;
   assign soundFileAmplitudes [6979] = 8'd135;
   assign soundFileAmplitudes [6980] = 8'd128;
   assign soundFileAmplitudes [6981] = 8'd119;
   assign soundFileAmplitudes [6982] = 8'd114;
   assign soundFileAmplitudes [6983] = 8'd128;
   assign soundFileAmplitudes [6984] = 8'd143;
   assign soundFileAmplitudes [6985] = 8'd127;
   assign soundFileAmplitudes [6986] = 8'd125;
   assign soundFileAmplitudes [6987] = 8'd123;
   assign soundFileAmplitudes [6988] = 8'd118;
   assign soundFileAmplitudes [6989] = 8'd97;
   assign soundFileAmplitudes [6990] = 8'd81;
   assign soundFileAmplitudes [6991] = 8'd90;
   assign soundFileAmplitudes [6992] = 8'd102;
   assign soundFileAmplitudes [6993] = 8'd110;
   assign soundFileAmplitudes [6994] = 8'd105;
   assign soundFileAmplitudes [6995] = 8'd102;
   assign soundFileAmplitudes [6996] = 8'd106;
   assign soundFileAmplitudes [6997] = 8'd113;
   assign soundFileAmplitudes [6998] = 8'd133;
   assign soundFileAmplitudes [6999] = 8'd152;
   assign soundFileAmplitudes [7000] = 8'd165;
   assign soundFileAmplitudes [7001] = 8'd176;
   assign soundFileAmplitudes [7002] = 8'd177;
   assign soundFileAmplitudes [7003] = 8'd169;
   assign soundFileAmplitudes [7004] = 8'd150;
   assign soundFileAmplitudes [7005] = 8'd143;
   assign soundFileAmplitudes [7006] = 8'd144;
   assign soundFileAmplitudes [7007] = 8'd138;
   assign soundFileAmplitudes [7008] = 8'd136;
   assign soundFileAmplitudes [7009] = 8'd129;
   assign soundFileAmplitudes [7010] = 8'd116;
   assign soundFileAmplitudes [7011] = 8'd100;
   assign soundFileAmplitudes [7012] = 8'd93;
   assign soundFileAmplitudes [7013] = 8'd105;
   assign soundFileAmplitudes [7014] = 8'd124;
   assign soundFileAmplitudes [7015] = 8'd134;
   assign soundFileAmplitudes [7016] = 8'd136;
   assign soundFileAmplitudes [7017] = 8'd129;
   assign soundFileAmplitudes [7018] = 8'd113;
   assign soundFileAmplitudes [7019] = 8'd116;
   assign soundFileAmplitudes [7020] = 8'd136;
   assign soundFileAmplitudes [7021] = 8'd143;
   assign soundFileAmplitudes [7022] = 8'd145;
   assign soundFileAmplitudes [7023] = 8'd148;
   assign soundFileAmplitudes [7024] = 8'd139;
   assign soundFileAmplitudes [7025] = 8'd125;
   assign soundFileAmplitudes [7026] = 8'd101;
   assign soundFileAmplitudes [7027] = 8'd88;
   assign soundFileAmplitudes [7028] = 8'd99;
   assign soundFileAmplitudes [7029] = 8'd110;
   assign soundFileAmplitudes [7030] = 8'd111;
   assign soundFileAmplitudes [7031] = 8'd100;
   assign soundFileAmplitudes [7032] = 8'd96;
   assign soundFileAmplitudes [7033] = 8'd99;
   assign soundFileAmplitudes [7034] = 8'd115;
   assign soundFileAmplitudes [7035] = 8'd138;
   assign soundFileAmplitudes [7036] = 8'd156;
   assign soundFileAmplitudes [7037] = 8'd167;
   assign soundFileAmplitudes [7038] = 8'd168;
   assign soundFileAmplitudes [7039] = 8'd171;
   assign soundFileAmplitudes [7040] = 8'd158;
   assign soundFileAmplitudes [7041] = 8'd138;
   assign soundFileAmplitudes [7042] = 8'd130;
   assign soundFileAmplitudes [7043] = 8'd122;
   assign soundFileAmplitudes [7044] = 8'd119;
   assign soundFileAmplitudes [7045] = 8'd117;
   assign soundFileAmplitudes [7046] = 8'd113;
   assign soundFileAmplitudes [7047] = 8'd104;
   assign soundFileAmplitudes [7048] = 8'd98;
   assign soundFileAmplitudes [7049] = 8'd101;
   assign soundFileAmplitudes [7050] = 8'd113;
   assign soundFileAmplitudes [7051] = 8'd127;
   assign soundFileAmplitudes [7052] = 8'd135;
   assign soundFileAmplitudes [7053] = 8'd136;
   assign soundFileAmplitudes [7054] = 8'd134;
   assign soundFileAmplitudes [7055] = 8'd125;
   assign soundFileAmplitudes [7056] = 8'd133;
   assign soundFileAmplitudes [7057] = 8'd143;
   assign soundFileAmplitudes [7058] = 8'd137;
   assign soundFileAmplitudes [7059] = 8'd130;
   assign soundFileAmplitudes [7060] = 8'd133;
   assign soundFileAmplitudes [7061] = 8'd137;
   assign soundFileAmplitudes [7062] = 8'd127;
   assign soundFileAmplitudes [7063] = 8'd104;
   assign soundFileAmplitudes [7064] = 8'd91;
   assign soundFileAmplitudes [7065] = 8'd100;
   assign soundFileAmplitudes [7066] = 8'd104;
   assign soundFileAmplitudes [7067] = 8'd106;
   assign soundFileAmplitudes [7068] = 8'd103;
   assign soundFileAmplitudes [7069] = 8'd102;
   assign soundFileAmplitudes [7070] = 8'd109;
   assign soundFileAmplitudes [7071] = 8'd122;
   assign soundFileAmplitudes [7072] = 8'd136;
   assign soundFileAmplitudes [7073] = 8'd155;
   assign soundFileAmplitudes [7074] = 8'd164;
   assign soundFileAmplitudes [7075] = 8'd168;
   assign soundFileAmplitudes [7076] = 8'd157;
   assign soundFileAmplitudes [7077] = 8'd143;
   assign soundFileAmplitudes [7078] = 8'd154;
   assign soundFileAmplitudes [7079] = 8'd157;
   assign soundFileAmplitudes [7080] = 8'd152;
   assign soundFileAmplitudes [7081] = 8'd133;
   assign soundFileAmplitudes [7082] = 8'd121;
   assign soundFileAmplitudes [7083] = 8'd104;
   assign soundFileAmplitudes [7084] = 8'd94;
   assign soundFileAmplitudes [7085] = 8'd97;
   assign soundFileAmplitudes [7086] = 8'd103;
   assign soundFileAmplitudes [7087] = 8'd124;
   assign soundFileAmplitudes [7088] = 8'd141;
   assign soundFileAmplitudes [7089] = 8'd141;
   assign soundFileAmplitudes [7090] = 8'd129;
   assign soundFileAmplitudes [7091] = 8'd118;
   assign soundFileAmplitudes [7092] = 8'd121;
   assign soundFileAmplitudes [7093] = 8'd141;
   assign soundFileAmplitudes [7094] = 8'd141;
   assign soundFileAmplitudes [7095] = 8'd141;
   assign soundFileAmplitudes [7096] = 8'd136;
   assign soundFileAmplitudes [7097] = 8'd128;
   assign soundFileAmplitudes [7098] = 8'd126;
   assign soundFileAmplitudes [7099] = 8'd98;
   assign soundFileAmplitudes [7100] = 8'd86;
   assign soundFileAmplitudes [7101] = 8'd97;
   assign soundFileAmplitudes [7102] = 8'd110;
   assign soundFileAmplitudes [7103] = 8'd120;
   assign soundFileAmplitudes [7104] = 8'd113;
   assign soundFileAmplitudes [7105] = 8'd109;
   assign soundFileAmplitudes [7106] = 8'd110;
   assign soundFileAmplitudes [7107] = 8'd114;
   assign soundFileAmplitudes [7108] = 8'd130;
   assign soundFileAmplitudes [7109] = 8'd145;
   assign soundFileAmplitudes [7110] = 8'd162;
   assign soundFileAmplitudes [7111] = 8'd173;
   assign soundFileAmplitudes [7112] = 8'd179;
   assign soundFileAmplitudes [7113] = 8'd165;
   assign soundFileAmplitudes [7114] = 8'd148;
   assign soundFileAmplitudes [7115] = 8'd145;
   assign soundFileAmplitudes [7116] = 8'd137;
   assign soundFileAmplitudes [7117] = 8'd128;
   assign soundFileAmplitudes [7118] = 8'd119;
   assign soundFileAmplitudes [7119] = 8'd117;
   assign soundFileAmplitudes [7120] = 8'd109;
   assign soundFileAmplitudes [7121] = 8'd96;
   assign soundFileAmplitudes [7122] = 8'd94;
   assign soundFileAmplitudes [7123] = 8'd104;
   assign soundFileAmplitudes [7124] = 8'd116;
   assign soundFileAmplitudes [7125] = 8'd127;
   assign soundFileAmplitudes [7126] = 8'd121;
   assign soundFileAmplitudes [7127] = 8'd116;
   assign soundFileAmplitudes [7128] = 8'd113;
   assign soundFileAmplitudes [7129] = 8'd108;
   assign soundFileAmplitudes [7130] = 8'd130;
   assign soundFileAmplitudes [7131] = 8'd151;
   assign soundFileAmplitudes [7132] = 8'd142;
   assign soundFileAmplitudes [7133] = 8'd135;
   assign soundFileAmplitudes [7134] = 8'd138;
   assign soundFileAmplitudes [7135] = 8'd139;
   assign soundFileAmplitudes [7136] = 8'd124;
   assign soundFileAmplitudes [7137] = 8'd105;
   assign soundFileAmplitudes [7138] = 8'd104;
   assign soundFileAmplitudes [7139] = 8'd111;
   assign soundFileAmplitudes [7140] = 8'd123;
   assign soundFileAmplitudes [7141] = 8'd120;
   assign soundFileAmplitudes [7142] = 8'd112;
   assign soundFileAmplitudes [7143] = 8'd114;
   assign soundFileAmplitudes [7144] = 8'd114;
   assign soundFileAmplitudes [7145] = 8'd130;
   assign soundFileAmplitudes [7146] = 8'd153;
   assign soundFileAmplitudes [7147] = 8'd163;
   assign soundFileAmplitudes [7148] = 8'd165;
   assign soundFileAmplitudes [7149] = 8'd153;
   assign soundFileAmplitudes [7150] = 8'd144;
   assign soundFileAmplitudes [7151] = 8'd141;
   assign soundFileAmplitudes [7152] = 8'd132;
   assign soundFileAmplitudes [7153] = 8'd125;
   assign soundFileAmplitudes [7154] = 8'd126;
   assign soundFileAmplitudes [7155] = 8'd123;
   assign soundFileAmplitudes [7156] = 8'd119;
   assign soundFileAmplitudes [7157] = 8'd108;
   assign soundFileAmplitudes [7158] = 8'd103;
   assign soundFileAmplitudes [7159] = 8'd104;
   assign soundFileAmplitudes [7160] = 8'd106;
   assign soundFileAmplitudes [7161] = 8'd111;
   assign soundFileAmplitudes [7162] = 8'd109;
   assign soundFileAmplitudes [7163] = 8'd115;
   assign soundFileAmplitudes [7164] = 8'd119;
   assign soundFileAmplitudes [7165] = 8'd123;
   assign soundFileAmplitudes [7166] = 8'd133;
   assign soundFileAmplitudes [7167] = 8'd148;
   assign soundFileAmplitudes [7168] = 8'd138;
   assign soundFileAmplitudes [7169] = 8'd132;
   assign soundFileAmplitudes [7170] = 8'd138;
   assign soundFileAmplitudes [7171] = 8'd144;
   assign soundFileAmplitudes [7172] = 8'd142;
   assign soundFileAmplitudes [7173] = 8'd109;
   assign soundFileAmplitudes [7174] = 8'd96;
   assign soundFileAmplitudes [7175] = 8'd102;
   assign soundFileAmplitudes [7176] = 8'd108;
   assign soundFileAmplitudes [7177] = 8'd112;
   assign soundFileAmplitudes [7178] = 8'd114;
   assign soundFileAmplitudes [7179] = 8'd113;
   assign soundFileAmplitudes [7180] = 8'd120;
   assign soundFileAmplitudes [7181] = 8'd132;
   assign soundFileAmplitudes [7182] = 8'd142;
   assign soundFileAmplitudes [7183] = 8'd146;
   assign soundFileAmplitudes [7184] = 8'd150;
   assign soundFileAmplitudes [7185] = 8'd149;
   assign soundFileAmplitudes [7186] = 8'd141;
   assign soundFileAmplitudes [7187] = 8'd145;
   assign soundFileAmplitudes [7188] = 8'd148;
   assign soundFileAmplitudes [7189] = 8'd154;
   assign soundFileAmplitudes [7190] = 8'd147;
   assign soundFileAmplitudes [7191] = 8'd140;
   assign soundFileAmplitudes [7192] = 8'd128;
   assign soundFileAmplitudes [7193] = 8'd119;
   assign soundFileAmplitudes [7194] = 8'd111;
   assign soundFileAmplitudes [7195] = 8'd104;
   assign soundFileAmplitudes [7196] = 8'd112;
   assign soundFileAmplitudes [7197] = 8'd120;
   assign soundFileAmplitudes [7198] = 8'd127;
   assign soundFileAmplitudes [7199] = 8'd114;
   assign soundFileAmplitudes [7200] = 8'd103;
   assign soundFileAmplitudes [7201] = 8'd99;
   assign soundFileAmplitudes [7202] = 8'd113;
   assign soundFileAmplitudes [7203] = 8'd133;
   assign soundFileAmplitudes [7204] = 8'd130;
   assign soundFileAmplitudes [7205] = 8'd127;
   assign soundFileAmplitudes [7206] = 8'd136;
   assign soundFileAmplitudes [7207] = 8'd136;
   assign soundFileAmplitudes [7208] = 8'd125;
   assign soundFileAmplitudes [7209] = 8'd97;
   assign soundFileAmplitudes [7210] = 8'd85;
   assign soundFileAmplitudes [7211] = 8'd98;
   assign soundFileAmplitudes [7212] = 8'd110;
   assign soundFileAmplitudes [7213] = 8'd130;
   assign soundFileAmplitudes [7214] = 8'd132;
   assign soundFileAmplitudes [7215] = 8'd123;
   assign soundFileAmplitudes [7216] = 8'd124;
   assign soundFileAmplitudes [7217] = 8'd133;
   assign soundFileAmplitudes [7218] = 8'd145;
   assign soundFileAmplitudes [7219] = 8'd155;
   assign soundFileAmplitudes [7220] = 8'd158;
   assign soundFileAmplitudes [7221] = 8'd160;
   assign soundFileAmplitudes [7222] = 8'd156;
   assign soundFileAmplitudes [7223] = 8'd149;
   assign soundFileAmplitudes [7224] = 8'd143;
   assign soundFileAmplitudes [7225] = 8'd146;
   assign soundFileAmplitudes [7226] = 8'd144;
   assign soundFileAmplitudes [7227] = 8'd138;
   assign soundFileAmplitudes [7228] = 8'd133;
   assign soundFileAmplitudes [7229] = 8'd121;
   assign soundFileAmplitudes [7230] = 8'd109;
   assign soundFileAmplitudes [7231] = 8'd101;
   assign soundFileAmplitudes [7232] = 8'd102;
   assign soundFileAmplitudes [7233] = 8'd111;
   assign soundFileAmplitudes [7234] = 8'd125;
   assign soundFileAmplitudes [7235] = 8'd123;
   assign soundFileAmplitudes [7236] = 8'd116;
   assign soundFileAmplitudes [7237] = 8'd112;
   assign soundFileAmplitudes [7238] = 8'd108;
   assign soundFileAmplitudes [7239] = 8'd110;
   assign soundFileAmplitudes [7240] = 8'd113;
   assign soundFileAmplitudes [7241] = 8'd113;
   assign soundFileAmplitudes [7242] = 8'd123;
   assign soundFileAmplitudes [7243] = 8'd133;
   assign soundFileAmplitudes [7244] = 8'd134;
   assign soundFileAmplitudes [7245] = 8'd114;
   assign soundFileAmplitudes [7246] = 8'd91;
   assign soundFileAmplitudes [7247] = 8'd96;
   assign soundFileAmplitudes [7248] = 8'd111;
   assign soundFileAmplitudes [7249] = 8'd129;
   assign soundFileAmplitudes [7250] = 8'd131;
   assign soundFileAmplitudes [7251] = 8'd133;
   assign soundFileAmplitudes [7252] = 8'd137;
   assign soundFileAmplitudes [7253] = 8'd147;
   assign soundFileAmplitudes [7254] = 8'd155;
   assign soundFileAmplitudes [7255] = 8'd155;
   assign soundFileAmplitudes [7256] = 8'd166;
   assign soundFileAmplitudes [7257] = 8'd163;
   assign soundFileAmplitudes [7258] = 8'd156;
   assign soundFileAmplitudes [7259] = 8'd152;
   assign soundFileAmplitudes [7260] = 8'd152;
   assign soundFileAmplitudes [7261] = 8'd146;
   assign soundFileAmplitudes [7262] = 8'd134;
   assign soundFileAmplitudes [7263] = 8'd134;
   assign soundFileAmplitudes [7264] = 8'd125;
   assign soundFileAmplitudes [7265] = 8'd114;
   assign soundFileAmplitudes [7266] = 8'd102;
   assign soundFileAmplitudes [7267] = 8'd101;
   assign soundFileAmplitudes [7268] = 8'd107;
   assign soundFileAmplitudes [7269] = 8'd116;
   assign soundFileAmplitudes [7270] = 8'd123;
   assign soundFileAmplitudes [7271] = 8'd116;
   assign soundFileAmplitudes [7272] = 8'd112;
   assign soundFileAmplitudes [7273] = 8'd109;
   assign soundFileAmplitudes [7274] = 8'd118;
   assign soundFileAmplitudes [7275] = 8'd128;
   assign soundFileAmplitudes [7276] = 8'd134;
   assign soundFileAmplitudes [7277] = 8'd127;
   assign soundFileAmplitudes [7278] = 8'd121;
   assign soundFileAmplitudes [7279] = 8'd122;
   assign soundFileAmplitudes [7280] = 8'd125;
   assign soundFileAmplitudes [7281] = 8'd120;
   assign soundFileAmplitudes [7282] = 8'd95;
   assign soundFileAmplitudes [7283] = 8'd78;
   assign soundFileAmplitudes [7284] = 8'd91;
   assign soundFileAmplitudes [7285] = 8'd116;
   assign soundFileAmplitudes [7286] = 8'd129;
   assign soundFileAmplitudes [7287] = 8'd125;
   assign soundFileAmplitudes [7288] = 8'd122;
   assign soundFileAmplitudes [7289] = 8'd129;
   assign soundFileAmplitudes [7290] = 8'd150;
   assign soundFileAmplitudes [7291] = 8'd165;
   assign soundFileAmplitudes [7292] = 8'd164;
   assign soundFileAmplitudes [7293] = 8'd166;
   assign soundFileAmplitudes [7294] = 8'd146;
   assign soundFileAmplitudes [7295] = 8'd143;
   assign soundFileAmplitudes [7296] = 8'd142;
   assign soundFileAmplitudes [7297] = 8'd134;
   assign soundFileAmplitudes [7298] = 8'd130;
   assign soundFileAmplitudes [7299] = 8'd120;
   assign soundFileAmplitudes [7300] = 8'd120;
   assign soundFileAmplitudes [7301] = 8'd112;
   assign soundFileAmplitudes [7302] = 8'd113;
   assign soundFileAmplitudes [7303] = 8'd119;
   assign soundFileAmplitudes [7304] = 8'd119;
   assign soundFileAmplitudes [7305] = 8'd125;
   assign soundFileAmplitudes [7306] = 8'd134;
   assign soundFileAmplitudes [7307] = 8'd136;
   assign soundFileAmplitudes [7308] = 8'd128;
   assign soundFileAmplitudes [7309] = 8'd117;
   assign soundFileAmplitudes [7310] = 8'd119;
   assign soundFileAmplitudes [7311] = 8'd126;
   assign soundFileAmplitudes [7312] = 8'd134;
   assign soundFileAmplitudes [7313] = 8'd133;
   assign soundFileAmplitudes [7314] = 8'd119;
   assign soundFileAmplitudes [7315] = 8'd114;
   assign soundFileAmplitudes [7316] = 8'd126;
   assign soundFileAmplitudes [7317] = 8'd127;
   assign soundFileAmplitudes [7318] = 8'd107;
   assign soundFileAmplitudes [7319] = 8'd72;
   assign soundFileAmplitudes [7320] = 8'd59;
   assign soundFileAmplitudes [7321] = 8'd78;
   assign soundFileAmplitudes [7322] = 8'd106;
   assign soundFileAmplitudes [7323] = 8'd128;
   assign soundFileAmplitudes [7324] = 8'd136;
   assign soundFileAmplitudes [7325] = 8'd143;
   assign soundFileAmplitudes [7326] = 8'd156;
   assign soundFileAmplitudes [7327] = 8'd165;
   assign soundFileAmplitudes [7328] = 8'd162;
   assign soundFileAmplitudes [7329] = 8'd159;
   assign soundFileAmplitudes [7330] = 8'd154;
   assign soundFileAmplitudes [7331] = 8'd154;
   assign soundFileAmplitudes [7332] = 8'd145;
   assign soundFileAmplitudes [7333] = 8'd143;
   assign soundFileAmplitudes [7334] = 8'd132;
   assign soundFileAmplitudes [7335] = 8'd127;
   assign soundFileAmplitudes [7336] = 8'd119;
   assign soundFileAmplitudes [7337] = 8'd116;
   assign soundFileAmplitudes [7338] = 8'd124;
   assign soundFileAmplitudes [7339] = 8'd123;
   assign soundFileAmplitudes [7340] = 8'd129;
   assign soundFileAmplitudes [7341] = 8'd126;
   assign soundFileAmplitudes [7342] = 8'd127;
   assign soundFileAmplitudes [7343] = 8'd121;
   assign soundFileAmplitudes [7344] = 8'd121;
   assign soundFileAmplitudes [7345] = 8'd118;
   assign soundFileAmplitudes [7346] = 8'd120;
   assign soundFileAmplitudes [7347] = 8'd125;
   assign soundFileAmplitudes [7348] = 8'd128;
   assign soundFileAmplitudes [7349] = 8'd127;
   assign soundFileAmplitudes [7350] = 8'd116;
   assign soundFileAmplitudes [7351] = 8'd104;
   assign soundFileAmplitudes [7352] = 8'd110;
   assign soundFileAmplitudes [7353] = 8'd113;
   assign soundFileAmplitudes [7354] = 8'd108;
   assign soundFileAmplitudes [7355] = 8'd99;
   assign soundFileAmplitudes [7356] = 8'd78;
   assign soundFileAmplitudes [7357] = 8'd86;
   assign soundFileAmplitudes [7358] = 8'd98;
   assign soundFileAmplitudes [7359] = 8'd114;
   assign soundFileAmplitudes [7360] = 8'd123;
   assign soundFileAmplitudes [7361] = 8'd135;
   assign soundFileAmplitudes [7362] = 8'd149;
   assign soundFileAmplitudes [7363] = 8'd164;
   assign soundFileAmplitudes [7364] = 8'd173;
   assign soundFileAmplitudes [7365] = 8'd169;
   assign soundFileAmplitudes [7366] = 8'd171;
   assign soundFileAmplitudes [7367] = 8'd161;
   assign soundFileAmplitudes [7368] = 8'd153;
   assign soundFileAmplitudes [7369] = 8'd147;
   assign soundFileAmplitudes [7370] = 8'd141;
   assign soundFileAmplitudes [7371] = 8'd138;
   assign soundFileAmplitudes [7372] = 8'd131;
   assign soundFileAmplitudes [7373] = 8'd134;
   assign soundFileAmplitudes [7374] = 8'd129;
   assign soundFileAmplitudes [7375] = 8'd124;
   assign soundFileAmplitudes [7376] = 8'd121;
   assign soundFileAmplitudes [7377] = 8'd113;
   assign soundFileAmplitudes [7378] = 8'd113;
   assign soundFileAmplitudes [7379] = 8'd118;
   assign soundFileAmplitudes [7380] = 8'd123;
   assign soundFileAmplitudes [7381] = 8'd127;
   assign soundFileAmplitudes [7382] = 8'd124;
   assign soundFileAmplitudes [7383] = 8'd122;
   assign soundFileAmplitudes [7384] = 8'd120;
   assign soundFileAmplitudes [7385] = 8'd109;
   assign soundFileAmplitudes [7386] = 8'd109;
   assign soundFileAmplitudes [7387] = 8'd111;
   assign soundFileAmplitudes [7388] = 8'd113;
   assign soundFileAmplitudes [7389] = 8'd117;
   assign soundFileAmplitudes [7390] = 8'd125;
   assign soundFileAmplitudes [7391] = 8'd122;
   assign soundFileAmplitudes [7392] = 8'd116;
   assign soundFileAmplitudes [7393] = 8'd102;
   assign soundFileAmplitudes [7394] = 8'd86;
   assign soundFileAmplitudes [7395] = 8'd96;
   assign soundFileAmplitudes [7396] = 8'd112;
   assign soundFileAmplitudes [7397] = 8'd134;
   assign soundFileAmplitudes [7398] = 8'd143;
   assign soundFileAmplitudes [7399] = 8'd145;
   assign soundFileAmplitudes [7400] = 8'd143;
   assign soundFileAmplitudes [7401] = 8'd139;
   assign soundFileAmplitudes [7402] = 8'd147;
   assign soundFileAmplitudes [7403] = 8'd155;
   assign soundFileAmplitudes [7404] = 8'd160;
   assign soundFileAmplitudes [7405] = 8'd160;
   assign soundFileAmplitudes [7406] = 8'd150;
   assign soundFileAmplitudes [7407] = 8'd138;
   assign soundFileAmplitudes [7408] = 8'd127;
   assign soundFileAmplitudes [7409] = 8'd127;
   assign soundFileAmplitudes [7410] = 8'd130;
   assign soundFileAmplitudes [7411] = 8'd131;
   assign soundFileAmplitudes [7412] = 8'd129;
   assign soundFileAmplitudes [7413] = 8'd115;
   assign soundFileAmplitudes [7414] = 8'd112;
   assign soundFileAmplitudes [7415] = 8'd113;
   assign soundFileAmplitudes [7416] = 8'd123;
   assign soundFileAmplitudes [7417] = 8'd131;
   assign soundFileAmplitudes [7418] = 8'd127;
   assign soundFileAmplitudes [7419] = 8'd129;
   assign soundFileAmplitudes [7420] = 8'd125;
   assign soundFileAmplitudes [7421] = 8'd126;
   assign soundFileAmplitudes [7422] = 8'd123;
   assign soundFileAmplitudes [7423] = 8'd112;
   assign soundFileAmplitudes [7424] = 8'd107;
   assign soundFileAmplitudes [7425] = 8'd106;
   assign soundFileAmplitudes [7426] = 8'd116;
   assign soundFileAmplitudes [7427] = 8'd131;
   assign soundFileAmplitudes [7428] = 8'd133;
   assign soundFileAmplitudes [7429] = 8'd126;
   assign soundFileAmplitudes [7430] = 8'd96;
   assign soundFileAmplitudes [7431] = 8'd85;
   assign soundFileAmplitudes [7432] = 8'd103;
   assign soundFileAmplitudes [7433] = 8'd120;
   assign soundFileAmplitudes [7434] = 8'd130;
   assign soundFileAmplitudes [7435] = 8'd131;
   assign soundFileAmplitudes [7436] = 8'd131;
   assign soundFileAmplitudes [7437] = 8'd136;
   assign soundFileAmplitudes [7438] = 8'd152;
   assign soundFileAmplitudes [7439] = 8'd150;
   assign soundFileAmplitudes [7440] = 8'd151;
   assign soundFileAmplitudes [7441] = 8'd147;
   assign soundFileAmplitudes [7442] = 8'd138;
   assign soundFileAmplitudes [7443] = 8'd132;
   assign soundFileAmplitudes [7444] = 8'd131;
   assign soundFileAmplitudes [7445] = 8'd131;
   assign soundFileAmplitudes [7446] = 8'd130;
   assign soundFileAmplitudes [7447] = 8'd134;
   assign soundFileAmplitudes [7448] = 8'd127;
   assign soundFileAmplitudes [7449] = 8'd118;
   assign soundFileAmplitudes [7450] = 8'd115;
   assign soundFileAmplitudes [7451] = 8'd116;
   assign soundFileAmplitudes [7452] = 8'd126;
   assign soundFileAmplitudes [7453] = 8'd138;
   assign soundFileAmplitudes [7454] = 8'd137;
   assign soundFileAmplitudes [7455] = 8'd136;
   assign soundFileAmplitudes [7456] = 8'd129;
   assign soundFileAmplitudes [7457] = 8'd118;
   assign soundFileAmplitudes [7458] = 8'd112;
   assign soundFileAmplitudes [7459] = 8'd109;
   assign soundFileAmplitudes [7460] = 8'd112;
   assign soundFileAmplitudes [7461] = 8'd112;
   assign soundFileAmplitudes [7462] = 8'd107;
   assign soundFileAmplitudes [7463] = 8'd116;
   assign soundFileAmplitudes [7464] = 8'd110;
   assign soundFileAmplitudes [7465] = 8'd104;
   assign soundFileAmplitudes [7466] = 8'd99;
   assign soundFileAmplitudes [7467] = 8'd87;
   assign soundFileAmplitudes [7468] = 8'd107;
   assign soundFileAmplitudes [7469] = 8'd130;
   assign soundFileAmplitudes [7470] = 8'd146;
   assign soundFileAmplitudes [7471] = 8'd145;
   assign soundFileAmplitudes [7472] = 8'd144;
   assign soundFileAmplitudes [7473] = 8'd143;
   assign soundFileAmplitudes [7474] = 8'd142;
   assign soundFileAmplitudes [7475] = 8'd149;
   assign soundFileAmplitudes [7476] = 8'd149;
   assign soundFileAmplitudes [7477] = 8'd151;
   assign soundFileAmplitudes [7478] = 8'd143;
   assign soundFileAmplitudes [7479] = 8'd141;
   assign soundFileAmplitudes [7480] = 8'd137;
   assign soundFileAmplitudes [7481] = 8'd130;
   assign soundFileAmplitudes [7482] = 8'd129;
   assign soundFileAmplitudes [7483] = 8'd123;
   assign soundFileAmplitudes [7484] = 8'd118;
   assign soundFileAmplitudes [7485] = 8'd106;
   assign soundFileAmplitudes [7486] = 8'd105;
   assign soundFileAmplitudes [7487] = 8'd114;
   assign soundFileAmplitudes [7488] = 8'd131;
   assign soundFileAmplitudes [7489] = 8'd144;
   assign soundFileAmplitudes [7490] = 8'd146;
   assign soundFileAmplitudes [7491] = 8'd136;
   assign soundFileAmplitudes [7492] = 8'd128;
   assign soundFileAmplitudes [7493] = 8'd128;
   assign soundFileAmplitudes [7494] = 8'd135;
   assign soundFileAmplitudes [7495] = 8'd135;
   assign soundFileAmplitudes [7496] = 8'd122;
   assign soundFileAmplitudes [7497] = 8'd122;
   assign soundFileAmplitudes [7498] = 8'd109;
   assign soundFileAmplitudes [7499] = 8'd109;
   assign soundFileAmplitudes [7500] = 8'd95;
   assign soundFileAmplitudes [7501] = 8'd82;
   assign soundFileAmplitudes [7502] = 8'd96;
   assign soundFileAmplitudes [7503] = 8'd114;
   assign soundFileAmplitudes [7504] = 8'd124;
   assign soundFileAmplitudes [7505] = 8'd123;
   assign soundFileAmplitudes [7506] = 8'd130;
   assign soundFileAmplitudes [7507] = 8'd137;
   assign soundFileAmplitudes [7508] = 8'd142;
   assign soundFileAmplitudes [7509] = 8'd151;
   assign soundFileAmplitudes [7510] = 8'd161;
   assign soundFileAmplitudes [7511] = 8'd164;
   assign soundFileAmplitudes [7512] = 8'd153;
   assign soundFileAmplitudes [7513] = 8'd133;
   assign soundFileAmplitudes [7514] = 8'd131;
   assign soundFileAmplitudes [7515] = 8'd135;
   assign soundFileAmplitudes [7516] = 8'd136;
   assign soundFileAmplitudes [7517] = 8'd134;
   assign soundFileAmplitudes [7518] = 8'd127;
   assign soundFileAmplitudes [7519] = 8'd114;
   assign soundFileAmplitudes [7520] = 8'd105;
   assign soundFileAmplitudes [7521] = 8'd104;
   assign soundFileAmplitudes [7522] = 8'd116;
   assign soundFileAmplitudes [7523] = 8'd130;
   assign soundFileAmplitudes [7524] = 8'd133;
   assign soundFileAmplitudes [7525] = 8'd132;
   assign soundFileAmplitudes [7526] = 8'd128;
   assign soundFileAmplitudes [7527] = 8'd125;
   assign soundFileAmplitudes [7528] = 8'd127;
   assign soundFileAmplitudes [7529] = 8'd128;
   assign soundFileAmplitudes [7530] = 8'd130;
   assign soundFileAmplitudes [7531] = 8'd129;
   assign soundFileAmplitudes [7532] = 8'd120;
   assign soundFileAmplitudes [7533] = 8'd117;
   assign soundFileAmplitudes [7534] = 8'd106;
   assign soundFileAmplitudes [7535] = 8'd103;
   assign soundFileAmplitudes [7536] = 8'd112;
   assign soundFileAmplitudes [7537] = 8'd119;
   assign soundFileAmplitudes [7538] = 8'd128;
   assign soundFileAmplitudes [7539] = 8'd130;
   assign soundFileAmplitudes [7540] = 8'd133;
   assign soundFileAmplitudes [7541] = 8'd134;
   assign soundFileAmplitudes [7542] = 8'd132;
   assign soundFileAmplitudes [7543] = 8'd135;
   assign soundFileAmplitudes [7544] = 8'd140;
   assign soundFileAmplitudes [7545] = 8'd143;
   assign soundFileAmplitudes [7546] = 8'd139;
   assign soundFileAmplitudes [7547] = 8'd131;
   assign soundFileAmplitudes [7548] = 8'd127;
   assign soundFileAmplitudes [7549] = 8'd125;
   assign soundFileAmplitudes [7550] = 8'd122;
   assign soundFileAmplitudes [7551] = 8'd124;
   assign soundFileAmplitudes [7552] = 8'd130;
   assign soundFileAmplitudes [7553] = 8'd123;
   assign soundFileAmplitudes [7554] = 8'd111;
   assign soundFileAmplitudes [7555] = 8'd108;
   assign soundFileAmplitudes [7556] = 8'd112;
   assign soundFileAmplitudes [7557] = 8'd118;
   assign soundFileAmplitudes [7558] = 8'd129;
   assign soundFileAmplitudes [7559] = 8'd136;
   assign soundFileAmplitudes [7560] = 8'd137;
   assign soundFileAmplitudes [7561] = 8'd137;
   assign soundFileAmplitudes [7562] = 8'd142;
   assign soundFileAmplitudes [7563] = 8'd143;
   assign soundFileAmplitudes [7564] = 8'd130;
   assign soundFileAmplitudes [7565] = 8'd121;
   assign soundFileAmplitudes [7566] = 8'd117;
   assign soundFileAmplitudes [7567] = 8'd120;
   assign soundFileAmplitudes [7568] = 8'd114;
   assign soundFileAmplitudes [7569] = 8'd107;
   assign soundFileAmplitudes [7570] = 8'd112;
   assign soundFileAmplitudes [7571] = 8'd116;
   assign soundFileAmplitudes [7572] = 8'd125;
   assign soundFileAmplitudes [7573] = 8'd126;
   assign soundFileAmplitudes [7574] = 8'd127;
   assign soundFileAmplitudes [7575] = 8'd132;
   assign soundFileAmplitudes [7576] = 8'd141;
   assign soundFileAmplitudes [7577] = 8'd152;
   assign soundFileAmplitudes [7578] = 8'd146;
   assign soundFileAmplitudes [7579] = 8'd146;
   assign soundFileAmplitudes [7580] = 8'd145;
   assign soundFileAmplitudes [7581] = 8'd139;
   assign soundFileAmplitudes [7582] = 8'd136;
   assign soundFileAmplitudes [7583] = 8'd126;
   assign soundFileAmplitudes [7584] = 8'd123;
   assign soundFileAmplitudes [7585] = 8'd119;
   assign soundFileAmplitudes [7586] = 8'd124;
   assign soundFileAmplitudes [7587] = 8'd113;
   assign soundFileAmplitudes [7588] = 8'd89;
   assign soundFileAmplitudes [7589] = 8'd85;
   assign soundFileAmplitudes [7590] = 8'd89;
   assign soundFileAmplitudes [7591] = 8'd107;
   assign soundFileAmplitudes [7592] = 8'd125;
   assign soundFileAmplitudes [7593] = 8'd136;
   assign soundFileAmplitudes [7594] = 8'd136;
   assign soundFileAmplitudes [7595] = 8'd133;
   assign soundFileAmplitudes [7596] = 8'd139;
   assign soundFileAmplitudes [7597] = 8'd138;
   assign soundFileAmplitudes [7598] = 8'd136;
   assign soundFileAmplitudes [7599] = 8'd144;
   assign soundFileAmplitudes [7600] = 8'd136;
   assign soundFileAmplitudes [7601] = 8'd131;
   assign soundFileAmplitudes [7602] = 8'd127;
   assign soundFileAmplitudes [7603] = 8'd112;
   assign soundFileAmplitudes [7604] = 8'd102;
   assign soundFileAmplitudes [7605] = 8'd93;
   assign soundFileAmplitudes [7606] = 8'd96;
   assign soundFileAmplitudes [7607] = 8'd104;
   assign soundFileAmplitudes [7608] = 8'd112;
   assign soundFileAmplitudes [7609] = 8'd124;
   assign soundFileAmplitudes [7610] = 8'd134;
   assign soundFileAmplitudes [7611] = 8'd139;
   assign soundFileAmplitudes [7612] = 8'd145;
   assign soundFileAmplitudes [7613] = 8'd149;
   assign soundFileAmplitudes [7614] = 8'd154;
   assign soundFileAmplitudes [7615] = 8'd153;
   assign soundFileAmplitudes [7616] = 8'd149;
   assign soundFileAmplitudes [7617] = 8'd139;
   assign soundFileAmplitudes [7618] = 8'd140;
   assign soundFileAmplitudes [7619] = 8'd152;
   assign soundFileAmplitudes [7620] = 8'd148;
   assign soundFileAmplitudes [7621] = 8'd144;
   assign soundFileAmplitudes [7622] = 8'd127;
   assign soundFileAmplitudes [7623] = 8'd107;
   assign soundFileAmplitudes [7624] = 8'd102;
   assign soundFileAmplitudes [7625] = 8'd102;
   assign soundFileAmplitudes [7626] = 8'd115;
   assign soundFileAmplitudes [7627] = 8'd126;
   assign soundFileAmplitudes [7628] = 8'd124;
   assign soundFileAmplitudes [7629] = 8'd116;
   assign soundFileAmplitudes [7630] = 8'd105;
   assign soundFileAmplitudes [7631] = 8'd109;
   assign soundFileAmplitudes [7632] = 8'd125;
   assign soundFileAmplitudes [7633] = 8'd134;
   assign soundFileAmplitudes [7634] = 8'd140;
   assign soundFileAmplitudes [7635] = 8'd142;
   assign soundFileAmplitudes [7636] = 8'd135;
   assign soundFileAmplitudes [7637] = 8'd130;
   assign soundFileAmplitudes [7638] = 8'd121;
   assign soundFileAmplitudes [7639] = 8'd106;
   assign soundFileAmplitudes [7640] = 8'd100;
   assign soundFileAmplitudes [7641] = 8'd111;
   assign soundFileAmplitudes [7642] = 8'd120;
   assign soundFileAmplitudes [7643] = 8'd122;
   assign soundFileAmplitudes [7644] = 8'd117;
   assign soundFileAmplitudes [7645] = 8'd109;
   assign soundFileAmplitudes [7646] = 8'd111;
   assign soundFileAmplitudes [7647] = 8'd126;
   assign soundFileAmplitudes [7648] = 8'd143;
   assign soundFileAmplitudes [7649] = 8'd151;
   assign soundFileAmplitudes [7650] = 8'd152;
   assign soundFileAmplitudes [7651] = 8'd150;
   assign soundFileAmplitudes [7652] = 8'd150;
   assign soundFileAmplitudes [7653] = 8'd151;
   assign soundFileAmplitudes [7654] = 8'd148;
   assign soundFileAmplitudes [7655] = 8'd151;
   assign soundFileAmplitudes [7656] = 8'd154;
   assign soundFileAmplitudes [7657] = 8'd143;
   assign soundFileAmplitudes [7658] = 8'd122;
   assign soundFileAmplitudes [7659] = 8'd108;
   assign soundFileAmplitudes [7660] = 8'd101;
   assign soundFileAmplitudes [7661] = 8'd112;
   assign soundFileAmplitudes [7662] = 8'd122;
   assign soundFileAmplitudes [7663] = 8'd120;
   assign soundFileAmplitudes [7664] = 8'd115;
   assign soundFileAmplitudes [7665] = 8'd111;
   assign soundFileAmplitudes [7666] = 8'd109;
   assign soundFileAmplitudes [7667] = 8'd111;
   assign soundFileAmplitudes [7668] = 8'd122;
   assign soundFileAmplitudes [7669] = 8'd113;
   assign soundFileAmplitudes [7670] = 8'd121;
   assign soundFileAmplitudes [7671] = 8'd124;
   assign soundFileAmplitudes [7672] = 8'd129;
   assign soundFileAmplitudes [7673] = 8'd130;
   assign soundFileAmplitudes [7674] = 8'd116;
   assign soundFileAmplitudes [7675] = 8'd123;
   assign soundFileAmplitudes [7676] = 8'd127;
   assign soundFileAmplitudes [7677] = 8'd134;
   assign soundFileAmplitudes [7678] = 8'd126;
   assign soundFileAmplitudes [7679] = 8'd121;
   assign soundFileAmplitudes [7680] = 8'd124;
   assign soundFileAmplitudes [7681] = 8'd132;
   assign soundFileAmplitudes [7682] = 8'd144;
   assign soundFileAmplitudes [7683] = 8'd151;
   assign soundFileAmplitudes [7684] = 8'd148;
   assign soundFileAmplitudes [7685] = 8'd143;
   assign soundFileAmplitudes [7686] = 8'd131;
   assign soundFileAmplitudes [7687] = 8'd130;
   assign soundFileAmplitudes [7688] = 8'd141;
   assign soundFileAmplitudes [7689] = 8'd142;
   assign soundFileAmplitudes [7690] = 8'd143;
   assign soundFileAmplitudes [7691] = 8'd139;
   assign soundFileAmplitudes [7692] = 8'd131;
   assign soundFileAmplitudes [7693] = 8'd110;
   assign soundFileAmplitudes [7694] = 8'd102;
   assign soundFileAmplitudes [7695] = 8'd111;
   assign soundFileAmplitudes [7696] = 8'd123;
   assign soundFileAmplitudes [7697] = 8'd136;
   assign soundFileAmplitudes [7698] = 8'd141;
   assign soundFileAmplitudes [7699] = 8'd130;
   assign soundFileAmplitudes [7700] = 8'd111;
   assign soundFileAmplitudes [7701] = 8'd105;
   assign soundFileAmplitudes [7702] = 8'd112;
   assign soundFileAmplitudes [7703] = 8'd122;
   assign soundFileAmplitudes [7704] = 8'd119;
   assign soundFileAmplitudes [7705] = 8'd125;
   assign soundFileAmplitudes [7706] = 8'd118;
   assign soundFileAmplitudes [7707] = 8'd116;
   assign soundFileAmplitudes [7708] = 8'd105;
   assign soundFileAmplitudes [7709] = 8'd97;
   assign soundFileAmplitudes [7710] = 8'd116;
   assign soundFileAmplitudes [7711] = 8'd128;
   assign soundFileAmplitudes [7712] = 8'd138;
   assign soundFileAmplitudes [7713] = 8'd133;
   assign soundFileAmplitudes [7714] = 8'd134;
   assign soundFileAmplitudes [7715] = 8'd130;
   assign soundFileAmplitudes [7716] = 8'd125;
   assign soundFileAmplitudes [7717] = 8'd127;
   assign soundFileAmplitudes [7718] = 8'd127;
   assign soundFileAmplitudes [7719] = 8'd129;
   assign soundFileAmplitudes [7720] = 8'd137;
   assign soundFileAmplitudes [7721] = 8'd135;
   assign soundFileAmplitudes [7722] = 8'd134;
   assign soundFileAmplitudes [7723] = 8'd140;
   assign soundFileAmplitudes [7724] = 8'd135;
   assign soundFileAmplitudes [7725] = 8'd124;
   assign soundFileAmplitudes [7726] = 8'd118;
   assign soundFileAmplitudes [7727] = 8'd119;
   assign soundFileAmplitudes [7728] = 8'd118;
   assign soundFileAmplitudes [7729] = 8'd116;
   assign soundFileAmplitudes [7730] = 8'd118;
   assign soundFileAmplitudes [7731] = 8'd127;
   assign soundFileAmplitudes [7732] = 8'd135;
   assign soundFileAmplitudes [7733] = 8'd139;
   assign soundFileAmplitudes [7734] = 8'd133;
   assign soundFileAmplitudes [7735] = 8'd128;
   assign soundFileAmplitudes [7736] = 8'd133;
   assign soundFileAmplitudes [7737] = 8'd133;
   assign soundFileAmplitudes [7738] = 8'd141;
   assign soundFileAmplitudes [7739] = 8'd129;
   assign soundFileAmplitudes [7740] = 8'd121;
   assign soundFileAmplitudes [7741] = 8'd129;
   assign soundFileAmplitudes [7742] = 8'd125;
   assign soundFileAmplitudes [7743] = 8'd126;
   assign soundFileAmplitudes [7744] = 8'd109;
   assign soundFileAmplitudes [7745] = 8'd104;
   assign soundFileAmplitudes [7746] = 8'd109;
   assign soundFileAmplitudes [7747] = 8'd111;
   assign soundFileAmplitudes [7748] = 8'd113;
   assign soundFileAmplitudes [7749] = 8'd122;
   assign soundFileAmplitudes [7750] = 8'd123;
   assign soundFileAmplitudes [7751] = 8'd117;
   assign soundFileAmplitudes [7752] = 8'd130;
   assign soundFileAmplitudes [7753] = 8'd136;
   assign soundFileAmplitudes [7754] = 8'd146;
   assign soundFileAmplitudes [7755] = 8'd144;
   assign soundFileAmplitudes [7756] = 8'd137;
   assign soundFileAmplitudes [7757] = 8'd139;
   assign soundFileAmplitudes [7758] = 8'd139;
   assign soundFileAmplitudes [7759] = 8'd132;
   assign soundFileAmplitudes [7760] = 8'd125;
   assign soundFileAmplitudes [7761] = 8'd123;
   assign soundFileAmplitudes [7762] = 8'd125;
   assign soundFileAmplitudes [7763] = 8'd114;
   assign soundFileAmplitudes [7764] = 8'd110;
   assign soundFileAmplitudes [7765] = 8'd117;
   assign soundFileAmplitudes [7766] = 8'd123;
   assign soundFileAmplitudes [7767] = 8'd129;
   assign soundFileAmplitudes [7768] = 8'd132;
   assign soundFileAmplitudes [7769] = 8'd132;
   assign soundFileAmplitudes [7770] = 8'd129;
   assign soundFileAmplitudes [7771] = 8'd135;
   assign soundFileAmplitudes [7772] = 8'd134;
   assign soundFileAmplitudes [7773] = 8'd147;
   assign soundFileAmplitudes [7774] = 8'd144;
   assign soundFileAmplitudes [7775] = 8'd144;
   assign soundFileAmplitudes [7776] = 8'd133;
   assign soundFileAmplitudes [7777] = 8'd125;
   assign soundFileAmplitudes [7778] = 8'd128;
   assign soundFileAmplitudes [7779] = 8'd101;
   assign soundFileAmplitudes [7780] = 8'd100;
   assign soundFileAmplitudes [7781] = 8'd103;
   assign soundFileAmplitudes [7782] = 8'd114;
   assign soundFileAmplitudes [7783] = 8'd131;
   assign soundFileAmplitudes [7784] = 8'd134;
   assign soundFileAmplitudes [7785] = 8'd131;
   assign soundFileAmplitudes [7786] = 8'd127;
   assign soundFileAmplitudes [7787] = 8'd123;
   assign soundFileAmplitudes [7788] = 8'd133;
   assign soundFileAmplitudes [7789] = 8'd139;
   assign soundFileAmplitudes [7790] = 8'd152;
   assign soundFileAmplitudes [7791] = 8'd149;
   assign soundFileAmplitudes [7792] = 8'd139;
   assign soundFileAmplitudes [7793] = 8'd138;
   assign soundFileAmplitudes [7794] = 8'd129;
   assign soundFileAmplitudes [7795] = 8'd124;
   assign soundFileAmplitudes [7796] = 8'd121;
   assign soundFileAmplitudes [7797] = 8'd120;
   assign soundFileAmplitudes [7798] = 8'd108;
   assign soundFileAmplitudes [7799] = 8'd104;
   assign soundFileAmplitudes [7800] = 8'd110;
   assign soundFileAmplitudes [7801] = 8'd109;
   assign soundFileAmplitudes [7802] = 8'd114;
   assign soundFileAmplitudes [7803] = 8'd123;
   assign soundFileAmplitudes [7804] = 8'd117;
   assign soundFileAmplitudes [7805] = 8'd112;
   assign soundFileAmplitudes [7806] = 8'd113;
   assign soundFileAmplitudes [7807] = 8'd117;
   assign soundFileAmplitudes [7808] = 8'd134;
   assign soundFileAmplitudes [7809] = 8'd137;
   assign soundFileAmplitudes [7810] = 8'd133;
   assign soundFileAmplitudes [7811] = 8'd142;
   assign soundFileAmplitudes [7812] = 8'd139;
   assign soundFileAmplitudes [7813] = 8'd144;
   assign soundFileAmplitudes [7814] = 8'd122;
   assign soundFileAmplitudes [7815] = 8'd113;
   assign soundFileAmplitudes [7816] = 8'd120;
   assign soundFileAmplitudes [7817] = 8'd132;
   assign soundFileAmplitudes [7818] = 8'd141;
   assign soundFileAmplitudes [7819] = 8'd129;
   assign soundFileAmplitudes [7820] = 8'd126;
   assign soundFileAmplitudes [7821] = 8'd120;
   assign soundFileAmplitudes [7822] = 8'd127;
   assign soundFileAmplitudes [7823] = 8'd136;
   assign soundFileAmplitudes [7824] = 8'd148;
   assign soundFileAmplitudes [7825] = 8'd160;
   assign soundFileAmplitudes [7826] = 8'd156;
   assign soundFileAmplitudes [7827] = 8'd143;
   assign soundFileAmplitudes [7828] = 8'd140;
   assign soundFileAmplitudes [7829] = 8'd144;
   assign soundFileAmplitudes [7830] = 8'd136;
   assign soundFileAmplitudes [7831] = 8'd130;
   assign soundFileAmplitudes [7832] = 8'd128;
   assign soundFileAmplitudes [7833] = 8'd120;
   assign soundFileAmplitudes [7834] = 8'd107;
   assign soundFileAmplitudes [7835] = 8'd94;
   assign soundFileAmplitudes [7836] = 8'd90;
   assign soundFileAmplitudes [7837] = 8'd100;
   assign soundFileAmplitudes [7838] = 8'd110;
   assign soundFileAmplitudes [7839] = 8'd109;
   assign soundFileAmplitudes [7840] = 8'd106;
   assign soundFileAmplitudes [7841] = 8'd110;
   assign soundFileAmplitudes [7842] = 8'd118;
   assign soundFileAmplitudes [7843] = 8'd121;
   assign soundFileAmplitudes [7844] = 8'd130;
   assign soundFileAmplitudes [7845] = 8'd127;
   assign soundFileAmplitudes [7846] = 8'd134;
   assign soundFileAmplitudes [7847] = 8'd136;
   assign soundFileAmplitudes [7848] = 8'd140;
   assign soundFileAmplitudes [7849] = 8'd137;
   assign soundFileAmplitudes [7850] = 8'd117;
   assign soundFileAmplitudes [7851] = 8'd119;
   assign soundFileAmplitudes [7852] = 8'd117;
   assign soundFileAmplitudes [7853] = 8'd124;
   assign soundFileAmplitudes [7854] = 8'd125;
   assign soundFileAmplitudes [7855] = 8'd122;
   assign soundFileAmplitudes [7856] = 8'd121;
   assign soundFileAmplitudes [7857] = 8'd124;
   assign soundFileAmplitudes [7858] = 8'd138;
   assign soundFileAmplitudes [7859] = 8'd146;
   assign soundFileAmplitudes [7860] = 8'd158;
   assign soundFileAmplitudes [7861] = 8'd159;
   assign soundFileAmplitudes [7862] = 8'd148;
   assign soundFileAmplitudes [7863] = 8'd140;
   assign soundFileAmplitudes [7864] = 8'd139;
   assign soundFileAmplitudes [7865] = 8'd138;
   assign soundFileAmplitudes [7866] = 8'd134;
   assign soundFileAmplitudes [7867] = 8'd133;
   assign soundFileAmplitudes [7868] = 8'd130;
   assign soundFileAmplitudes [7869] = 8'd112;
   assign soundFileAmplitudes [7870] = 8'd95;
   assign soundFileAmplitudes [7871] = 8'd91;
   assign soundFileAmplitudes [7872] = 8'd88;
   assign soundFileAmplitudes [7873] = 8'd99;
   assign soundFileAmplitudes [7874] = 8'd113;
   assign soundFileAmplitudes [7875] = 8'd116;
   assign soundFileAmplitudes [7876] = 8'd116;
   assign soundFileAmplitudes [7877] = 8'd112;
   assign soundFileAmplitudes [7878] = 8'd115;
   assign soundFileAmplitudes [7879] = 8'd126;
   assign soundFileAmplitudes [7880] = 8'd135;
   assign soundFileAmplitudes [7881] = 8'd141;
   assign soundFileAmplitudes [7882] = 8'd144;
   assign soundFileAmplitudes [7883] = 8'd134;
   assign soundFileAmplitudes [7884] = 8'd134;
   assign soundFileAmplitudes [7885] = 8'd120;
   assign soundFileAmplitudes [7886] = 8'd103;
   assign soundFileAmplitudes [7887] = 8'd109;
   assign soundFileAmplitudes [7888] = 8'd116;
   assign soundFileAmplitudes [7889] = 8'd126;
   assign soundFileAmplitudes [7890] = 8'd128;
   assign soundFileAmplitudes [7891] = 8'd130;
   assign soundFileAmplitudes [7892] = 8'd132;
   assign soundFileAmplitudes [7893] = 8'd143;
   assign soundFileAmplitudes [7894] = 8'd156;
   assign soundFileAmplitudes [7895] = 8'd162;
   assign soundFileAmplitudes [7896] = 8'd163;
   assign soundFileAmplitudes [7897] = 8'd149;
   assign soundFileAmplitudes [7898] = 8'd146;
   assign soundFileAmplitudes [7899] = 8'd152;
   assign soundFileAmplitudes [7900] = 8'd149;
   assign soundFileAmplitudes [7901] = 8'd142;
   assign soundFileAmplitudes [7902] = 8'd136;
   assign soundFileAmplitudes [7903] = 8'd132;
   assign soundFileAmplitudes [7904] = 8'd116;
   assign soundFileAmplitudes [7905] = 8'd96;
   assign soundFileAmplitudes [7906] = 8'd90;
   assign soundFileAmplitudes [7907] = 8'd94;
   assign soundFileAmplitudes [7908] = 8'd104;
   assign soundFileAmplitudes [7909] = 8'd111;
   assign soundFileAmplitudes [7910] = 8'd111;
   assign soundFileAmplitudes [7911] = 8'd110;
   assign soundFileAmplitudes [7912] = 8'd113;
   assign soundFileAmplitudes [7913] = 8'd117;
   assign soundFileAmplitudes [7914] = 8'd125;
   assign soundFileAmplitudes [7915] = 8'd130;
   assign soundFileAmplitudes [7916] = 8'd133;
   assign soundFileAmplitudes [7917] = 8'd129;
   assign soundFileAmplitudes [7918] = 8'd135;
   assign soundFileAmplitudes [7919] = 8'd134;
   assign soundFileAmplitudes [7920] = 8'd122;
   assign soundFileAmplitudes [7921] = 8'd112;
   assign soundFileAmplitudes [7922] = 8'd101;
   assign soundFileAmplitudes [7923] = 8'd101;
   assign soundFileAmplitudes [7924] = 8'd104;
   assign soundFileAmplitudes [7925] = 8'd121;
   assign soundFileAmplitudes [7926] = 8'd132;
   assign soundFileAmplitudes [7927] = 8'd138;
   assign soundFileAmplitudes [7928] = 8'd137;
   assign soundFileAmplitudes [7929] = 8'd137;
   assign soundFileAmplitudes [7930] = 8'd141;
   assign soundFileAmplitudes [7931] = 8'd149;
   assign soundFileAmplitudes [7932] = 8'd172;
   assign soundFileAmplitudes [7933] = 8'd169;
   assign soundFileAmplitudes [7934] = 8'd160;
   assign soundFileAmplitudes [7935] = 8'd154;
   assign soundFileAmplitudes [7936] = 8'd141;
   assign soundFileAmplitudes [7937] = 8'd136;
   assign soundFileAmplitudes [7938] = 8'd132;
   assign soundFileAmplitudes [7939] = 8'd122;
   assign soundFileAmplitudes [7940] = 8'd108;
   assign soundFileAmplitudes [7941] = 8'd102;
   assign soundFileAmplitudes [7942] = 8'd107;
   assign soundFileAmplitudes [7943] = 8'd112;
   assign soundFileAmplitudes [7944] = 8'd116;
   assign soundFileAmplitudes [7945] = 8'd114;
   assign soundFileAmplitudes [7946] = 8'd109;
   assign soundFileAmplitudes [7947] = 8'd112;
   assign soundFileAmplitudes [7948] = 8'd124;
   assign soundFileAmplitudes [7949] = 8'd130;
   assign soundFileAmplitudes [7950] = 8'd141;
   assign soundFileAmplitudes [7951] = 8'd138;
   assign soundFileAmplitudes [7952] = 8'd127;
   assign soundFileAmplitudes [7953] = 8'd129;
   assign soundFileAmplitudes [7954] = 8'd132;
   assign soundFileAmplitudes [7955] = 8'd136;
   assign soundFileAmplitudes [7956] = 8'd113;
   assign soundFileAmplitudes [7957] = 8'd108;
   assign soundFileAmplitudes [7958] = 8'd124;
   assign soundFileAmplitudes [7959] = 8'd132;
   assign soundFileAmplitudes [7960] = 8'd126;
   assign soundFileAmplitudes [7961] = 8'd111;
   assign soundFileAmplitudes [7962] = 8'd100;
   assign soundFileAmplitudes [7963] = 8'd105;
   assign soundFileAmplitudes [7964] = 8'd127;
   assign soundFileAmplitudes [7965] = 8'd145;
   assign soundFileAmplitudes [7966] = 8'd154;
   assign soundFileAmplitudes [7967] = 8'd151;
   assign soundFileAmplitudes [7968] = 8'd146;
   assign soundFileAmplitudes [7969] = 8'd138;
   assign soundFileAmplitudes [7970] = 8'd152;
   assign soundFileAmplitudes [7971] = 8'd150;
   assign soundFileAmplitudes [7972] = 8'd138;
   assign soundFileAmplitudes [7973] = 8'd129;
   assign soundFileAmplitudes [7974] = 8'd123;
   assign soundFileAmplitudes [7975] = 8'd124;
   assign soundFileAmplitudes [7976] = 8'd114;
   assign soundFileAmplitudes [7977] = 8'd105;
   assign soundFileAmplitudes [7978] = 8'd95;
   assign soundFileAmplitudes [7979] = 8'd99;
   assign soundFileAmplitudes [7980] = 8'd110;
   assign soundFileAmplitudes [7981] = 8'd118;
   assign soundFileAmplitudes [7982] = 8'd121;
   assign soundFileAmplitudes [7983] = 8'd121;
   assign soundFileAmplitudes [7984] = 8'd124;
   assign soundFileAmplitudes [7985] = 8'd129;
   assign soundFileAmplitudes [7986] = 8'd140;
   assign soundFileAmplitudes [7987] = 8'd138;
   assign soundFileAmplitudes [7988] = 8'd133;
   assign soundFileAmplitudes [7989] = 8'd133;
   assign soundFileAmplitudes [7990] = 8'd131;
   assign soundFileAmplitudes [7991] = 8'd133;
   assign soundFileAmplitudes [7992] = 8'd117;
   assign soundFileAmplitudes [7993] = 8'd105;
   assign soundFileAmplitudes [7994] = 8'd111;
   assign soundFileAmplitudes [7995] = 8'd114;
   assign soundFileAmplitudes [7996] = 8'd116;
   assign soundFileAmplitudes [7997] = 8'd121;
   assign soundFileAmplitudes [7998] = 8'd118;
   assign soundFileAmplitudes [7999] = 8'd112;
   assign soundFileAmplitudes [8000] = 8'd114;
   assign soundFileAmplitudes [8001] = 8'd123;
   assign soundFileAmplitudes [8002] = 8'd138;
   assign soundFileAmplitudes [8003] = 8'd149;
   assign soundFileAmplitudes [8004] = 8'd150;
   assign soundFileAmplitudes [8005] = 8'd145;
   assign soundFileAmplitudes [8006] = 8'd131;
   assign soundFileAmplitudes [8007] = 8'd121;
   assign soundFileAmplitudes [8008] = 8'd127;
   assign soundFileAmplitudes [8009] = 8'd136;
   assign soundFileAmplitudes [8010] = 8'd150;
   assign soundFileAmplitudes [8011] = 8'd149;
   assign soundFileAmplitudes [8012] = 8'd141;
   assign soundFileAmplitudes [8013] = 8'd139;
   assign soundFileAmplitudes [8014] = 8'd131;
   assign soundFileAmplitudes [8015] = 8'd121;
   assign soundFileAmplitudes [8016] = 8'd125;
   assign soundFileAmplitudes [8017] = 8'd134;
   assign soundFileAmplitudes [8018] = 8'd136;
   assign soundFileAmplitudes [8019] = 8'd132;
   assign soundFileAmplitudes [8020] = 8'd120;
   assign soundFileAmplitudes [8021] = 8'd114;
   assign soundFileAmplitudes [8022] = 8'd117;
   assign soundFileAmplitudes [8023] = 8'd121;
   assign soundFileAmplitudes [8024] = 8'd126;
   assign soundFileAmplitudes [8025] = 8'd129;
   assign soundFileAmplitudes [8026] = 8'd136;
   assign soundFileAmplitudes [8027] = 8'd138;
   assign soundFileAmplitudes [8028] = 8'd132;
   assign soundFileAmplitudes [8029] = 8'd126;
   assign soundFileAmplitudes [8030] = 8'd123;
   assign soundFileAmplitudes [8031] = 8'd124;
   assign soundFileAmplitudes [8032] = 8'd130;
   assign soundFileAmplitudes [8033] = 8'd126;
   assign soundFileAmplitudes [8034] = 8'd117;
   assign soundFileAmplitudes [8035] = 8'd113;
   assign soundFileAmplitudes [8036] = 8'd108;
   assign soundFileAmplitudes [8037] = 8'd108;
   assign soundFileAmplitudes [8038] = 8'd118;
   assign soundFileAmplitudes [8039] = 8'd123;
   assign soundFileAmplitudes [8040] = 8'd127;
   assign soundFileAmplitudes [8041] = 8'd127;
   assign soundFileAmplitudes [8042] = 8'd131;
   assign soundFileAmplitudes [8043] = 8'd131;
   assign soundFileAmplitudes [8044] = 8'd125;
   assign soundFileAmplitudes [8045] = 8'd139;
   assign soundFileAmplitudes [8046] = 8'd142;
   assign soundFileAmplitudes [8047] = 8'd146;
   assign soundFileAmplitudes [8048] = 8'd151;
   assign soundFileAmplitudes [8049] = 8'd154;
   assign soundFileAmplitudes [8050] = 8'd151;
   assign soundFileAmplitudes [8051] = 8'd138;
   assign soundFileAmplitudes [8052] = 8'd131;
   assign soundFileAmplitudes [8053] = 8'd130;
   assign soundFileAmplitudes [8054] = 8'd128;
   assign soundFileAmplitudes [8055] = 8'd124;
   assign soundFileAmplitudes [8056] = 8'd119;
   assign soundFileAmplitudes [8057] = 8'd117;
   assign soundFileAmplitudes [8058] = 8'd112;
   assign soundFileAmplitudes [8059] = 8'd104;
   assign soundFileAmplitudes [8060] = 8'd103;
   assign soundFileAmplitudes [8061] = 8'd110;
   assign soundFileAmplitudes [8062] = 8'd121;
   assign soundFileAmplitudes [8063] = 8'd131;
   assign soundFileAmplitudes [8064] = 8'd134;
   assign soundFileAmplitudes [8065] = 8'd125;
   assign soundFileAmplitudes [8066] = 8'd122;
   assign soundFileAmplitudes [8067] = 8'd127;
   assign soundFileAmplitudes [8068] = 8'd136;
   assign soundFileAmplitudes [8069] = 8'd128;
   assign soundFileAmplitudes [8070] = 8'd126;
   assign soundFileAmplitudes [8071] = 8'd118;
   assign soundFileAmplitudes [8072] = 8'd108;
   assign soundFileAmplitudes [8073] = 8'd102;
   assign soundFileAmplitudes [8074] = 8'd101;
   assign soundFileAmplitudes [8075] = 8'd114;
   assign soundFileAmplitudes [8076] = 8'd120;
   assign soundFileAmplitudes [8077] = 8'd129;
   assign soundFileAmplitudes [8078] = 8'd125;
   assign soundFileAmplitudes [8079] = 8'd123;
   assign soundFileAmplitudes [8080] = 8'd133;
   assign soundFileAmplitudes [8081] = 8'd146;
   assign soundFileAmplitudes [8082] = 8'd154;
   assign soundFileAmplitudes [8083] = 8'd155;
   assign soundFileAmplitudes [8084] = 8'd156;
   assign soundFileAmplitudes [8085] = 8'd153;
   assign soundFileAmplitudes [8086] = 8'd140;
   assign soundFileAmplitudes [8087] = 8'd132;
   assign soundFileAmplitudes [8088] = 8'd134;
   assign soundFileAmplitudes [8089] = 8'd133;
   assign soundFileAmplitudes [8090] = 8'd126;
   assign soundFileAmplitudes [8091] = 8'd116;
   assign soundFileAmplitudes [8092] = 8'd109;
   assign soundFileAmplitudes [8093] = 8'd106;
   assign soundFileAmplitudes [8094] = 8'd100;
   assign soundFileAmplitudes [8095] = 8'd101;
   assign soundFileAmplitudes [8096] = 8'd109;
   assign soundFileAmplitudes [8097] = 8'd113;
   assign soundFileAmplitudes [8098] = 8'd116;
   assign soundFileAmplitudes [8099] = 8'd120;
   assign soundFileAmplitudes [8100] = 8'd126;
   assign soundFileAmplitudes [8101] = 8'd133;
   assign soundFileAmplitudes [8102] = 8'd134;
   assign soundFileAmplitudes [8103] = 8'd133;
   assign soundFileAmplitudes [8104] = 8'd136;
   assign soundFileAmplitudes [8105] = 8'd132;
   assign soundFileAmplitudes [8106] = 8'd129;
   assign soundFileAmplitudes [8107] = 8'd115;
   assign soundFileAmplitudes [8108] = 8'd115;
   assign soundFileAmplitudes [8109] = 8'd116;
   assign soundFileAmplitudes [8110] = 8'd117;
   assign soundFileAmplitudes [8111] = 8'd125;
   assign soundFileAmplitudes [8112] = 8'd124;
   assign soundFileAmplitudes [8113] = 8'd128;
   assign soundFileAmplitudes [8114] = 8'd125;
   assign soundFileAmplitudes [8115] = 8'd129;
   assign soundFileAmplitudes [8116] = 8'd139;
   assign soundFileAmplitudes [8117] = 8'd146;
   assign soundFileAmplitudes [8118] = 8'd146;
   assign soundFileAmplitudes [8119] = 8'd144;
   assign soundFileAmplitudes [8120] = 8'd141;
   assign soundFileAmplitudes [8121] = 8'd136;
   assign soundFileAmplitudes [8122] = 8'd130;
   assign soundFileAmplitudes [8123] = 8'd129;
   assign soundFileAmplitudes [8124] = 8'd131;
   assign soundFileAmplitudes [8125] = 8'd126;
   assign soundFileAmplitudes [8126] = 8'd114;
   assign soundFileAmplitudes [8127] = 8'd101;
   assign soundFileAmplitudes [8128] = 8'd107;
   assign soundFileAmplitudes [8129] = 8'd115;
   assign soundFileAmplitudes [8130] = 8'd117;
   assign soundFileAmplitudes [8131] = 8'd121;
   assign soundFileAmplitudes [8132] = 8'd113;
   assign soundFileAmplitudes [8133] = 8'd115;
   assign soundFileAmplitudes [8134] = 8'd135;
   assign soundFileAmplitudes [8135] = 8'd141;
   assign soundFileAmplitudes [8136] = 8'd137;
   assign soundFileAmplitudes [8137] = 8'd135;
   assign soundFileAmplitudes [8138] = 8'd134;
   assign soundFileAmplitudes [8139] = 8'd139;
   assign soundFileAmplitudes [8140] = 8'd136;
   assign soundFileAmplitudes [8141] = 8'd113;
   assign soundFileAmplitudes [8142] = 8'd100;
   assign soundFileAmplitudes [8143] = 8'd103;
   assign soundFileAmplitudes [8144] = 8'd113;
   assign soundFileAmplitudes [8145] = 8'd124;
   assign soundFileAmplitudes [8146] = 8'd130;
   assign soundFileAmplitudes [8147] = 8'd132;
   assign soundFileAmplitudes [8148] = 8'd133;
   assign soundFileAmplitudes [8149] = 8'd132;
   assign soundFileAmplitudes [8150] = 8'd132;
   assign soundFileAmplitudes [8151] = 8'd143;
   assign soundFileAmplitudes [8152] = 8'd154;
   assign soundFileAmplitudes [8153] = 8'd156;
   assign soundFileAmplitudes [8154] = 8'd152;
   assign soundFileAmplitudes [8155] = 8'd146;
   assign soundFileAmplitudes [8156] = 8'd145;
   assign soundFileAmplitudes [8157] = 8'd135;
   assign soundFileAmplitudes [8158] = 8'd122;
   assign soundFileAmplitudes [8159] = 8'd120;
   assign soundFileAmplitudes [8160] = 8'd110;
   assign soundFileAmplitudes [8161] = 8'd111;
   assign soundFileAmplitudes [8162] = 8'd114;
   assign soundFileAmplitudes [8163] = 8'd117;
   assign soundFileAmplitudes [8164] = 8'd120;
   assign soundFileAmplitudes [8165] = 8'd102;
   assign soundFileAmplitudes [8166] = 8'd104;
   assign soundFileAmplitudes [8167] = 8'd117;
   assign soundFileAmplitudes [8168] = 8'd131;
   assign soundFileAmplitudes [8169] = 8'd147;
   assign soundFileAmplitudes [8170] = 8'd141;
   assign soundFileAmplitudes [8171] = 8'd134;
   assign soundFileAmplitudes [8172] = 8'd129;
   assign soundFileAmplitudes [8173] = 8'd125;
   assign soundFileAmplitudes [8174] = 8'd126;
   assign soundFileAmplitudes [8175] = 8'd119;
   assign soundFileAmplitudes [8176] = 8'd111;
   assign soundFileAmplitudes [8177] = 8'd111;
   assign soundFileAmplitudes [8178] = 8'd113;
   assign soundFileAmplitudes [8179] = 8'd109;
   assign soundFileAmplitudes [8180] = 8'd113;
   assign soundFileAmplitudes [8181] = 8'd133;
   assign soundFileAmplitudes [8182] = 8'd139;
   assign soundFileAmplitudes [8183] = 8'd145;
   assign soundFileAmplitudes [8184] = 8'd140;
   assign soundFileAmplitudes [8185] = 8'd132;
   assign soundFileAmplitudes [8186] = 8'd143;
   assign soundFileAmplitudes [8187] = 8'd153;
   assign soundFileAmplitudes [8188] = 8'd161;
   assign soundFileAmplitudes [8189] = 8'd157;
   assign soundFileAmplitudes [8190] = 8'd145;
   assign soundFileAmplitudes [8191] = 8'd137;
   assign soundFileAmplitudes [8192] = 8'd121;
   assign soundFileAmplitudes [8193] = 8'd110;
   assign soundFileAmplitudes [8194] = 8'd111;
   assign soundFileAmplitudes [8195] = 8'd110;
   assign soundFileAmplitudes [8196] = 8'd111;
   assign soundFileAmplitudes [8197] = 8'd107;
   assign soundFileAmplitudes [8198] = 8'd104;
   assign soundFileAmplitudes [8199] = 8'd112;
   assign soundFileAmplitudes [8200] = 8'd116;
   assign soundFileAmplitudes [8201] = 8'd118;
   assign soundFileAmplitudes [8202] = 8'd121;
   assign soundFileAmplitudes [8203] = 8'd125;
   assign soundFileAmplitudes [8204] = 8'd128;
   assign soundFileAmplitudes [8205] = 8'd128;
   assign soundFileAmplitudes [8206] = 8'd130;
   assign soundFileAmplitudes [8207] = 8'd125;
   assign soundFileAmplitudes [8208] = 8'd123;
   assign soundFileAmplitudes [8209] = 8'd122;
   assign soundFileAmplitudes [8210] = 8'd114;
   assign soundFileAmplitudes [8211] = 8'd117;
   assign soundFileAmplitudes [8212] = 8'd122;
   assign soundFileAmplitudes [8213] = 8'd116;
   assign soundFileAmplitudes [8214] = 8'd119;
   assign soundFileAmplitudes [8215] = 8'd126;
   assign soundFileAmplitudes [8216] = 8'd127;
   assign soundFileAmplitudes [8217] = 8'd135;
   assign soundFileAmplitudes [8218] = 8'd138;
   assign soundFileAmplitudes [8219] = 8'd144;
   assign soundFileAmplitudes [8220] = 8'd145;
   assign soundFileAmplitudes [8221] = 8'd153;
   assign soundFileAmplitudes [8222] = 8'd159;
   assign soundFileAmplitudes [8223] = 8'd158;
   assign soundFileAmplitudes [8224] = 8'd150;
   assign soundFileAmplitudes [8225] = 8'd130;
   assign soundFileAmplitudes [8226] = 8'd123;
   assign soundFileAmplitudes [8227] = 8'd115;
   assign soundFileAmplitudes [8228] = 8'd103;
   assign soundFileAmplitudes [8229] = 8'd103;
   assign soundFileAmplitudes [8230] = 8'd107;
   assign soundFileAmplitudes [8231] = 8'd108;
   assign soundFileAmplitudes [8232] = 8'd110;
   assign soundFileAmplitudes [8233] = 8'd108;
   assign soundFileAmplitudes [8234] = 8'd117;
   assign soundFileAmplitudes [8235] = 8'd126;
   assign soundFileAmplitudes [8236] = 8'd136;
   assign soundFileAmplitudes [8237] = 8'd141;
   assign soundFileAmplitudes [8238] = 8'd130;
   assign soundFileAmplitudes [8239] = 8'd134;
   assign soundFileAmplitudes [8240] = 8'd145;
   assign soundFileAmplitudes [8241] = 8'd143;
   assign soundFileAmplitudes [8242] = 8'd123;
   assign soundFileAmplitudes [8243] = 8'd110;
   assign soundFileAmplitudes [8244] = 8'd111;
   assign soundFileAmplitudes [8245] = 8'd123;
   assign soundFileAmplitudes [8246] = 8'd123;
   assign soundFileAmplitudes [8247] = 8'd119;
   assign soundFileAmplitudes [8248] = 8'd107;
   assign soundFileAmplitudes [8249] = 8'd98;
   assign soundFileAmplitudes [8250] = 8'd108;
   assign soundFileAmplitudes [8251] = 8'd123;
   assign soundFileAmplitudes [8252] = 8'd134;
   assign soundFileAmplitudes [8253] = 8'd143;
   assign soundFileAmplitudes [8254] = 8'd150;
   assign soundFileAmplitudes [8255] = 8'd150;
   assign soundFileAmplitudes [8256] = 8'd147;
   assign soundFileAmplitudes [8257] = 8'd143;
   assign soundFileAmplitudes [8258] = 8'd141;
   assign soundFileAmplitudes [8259] = 8'd141;
   assign soundFileAmplitudes [8260] = 8'd134;
   assign soundFileAmplitudes [8261] = 8'd127;
   assign soundFileAmplitudes [8262] = 8'd117;
   assign soundFileAmplitudes [8263] = 8'd99;
   assign soundFileAmplitudes [8264] = 8'd106;
   assign soundFileAmplitudes [8265] = 8'd116;
   assign soundFileAmplitudes [8266] = 8'd116;
   assign soundFileAmplitudes [8267] = 8'd118;
   assign soundFileAmplitudes [8268] = 8'd118;
   assign soundFileAmplitudes [8269] = 8'd122;
   assign soundFileAmplitudes [8270] = 8'd129;
   assign soundFileAmplitudes [8271] = 8'd117;
   assign soundFileAmplitudes [8272] = 8'd118;
   assign soundFileAmplitudes [8273] = 8'd123;
   assign soundFileAmplitudes [8274] = 8'd129;
   assign soundFileAmplitudes [8275] = 8'd135;
   assign soundFileAmplitudes [8276] = 8'd123;
   assign soundFileAmplitudes [8277] = 8'd126;
   assign soundFileAmplitudes [8278] = 8'd126;
   assign soundFileAmplitudes [8279] = 8'd133;
   assign soundFileAmplitudes [8280] = 8'd133;
   assign soundFileAmplitudes [8281] = 8'd130;
   assign soundFileAmplitudes [8282] = 8'd129;
   assign soundFileAmplitudes [8283] = 8'd126;
   assign soundFileAmplitudes [8284] = 8'd122;
   assign soundFileAmplitudes [8285] = 8'd122;
   assign soundFileAmplitudes [8286] = 8'd124;
   assign soundFileAmplitudes [8287] = 8'd136;
   assign soundFileAmplitudes [8288] = 8'd146;
   assign soundFileAmplitudes [8289] = 8'd141;
   assign soundFileAmplitudes [8290] = 8'd140;
   assign soundFileAmplitudes [8291] = 8'd127;
   assign soundFileAmplitudes [8292] = 8'd117;
   assign soundFileAmplitudes [8293] = 8'd126;
   assign soundFileAmplitudes [8294] = 8'd131;
   assign soundFileAmplitudes [8295] = 8'd127;
   assign soundFileAmplitudes [8296] = 8'd132;
   assign soundFileAmplitudes [8297] = 8'd132;
   assign soundFileAmplitudes [8298] = 8'd128;
   assign soundFileAmplitudes [8299] = 8'd114;
   assign soundFileAmplitudes [8300] = 8'd109;
   assign soundFileAmplitudes [8301] = 8'd118;
   assign soundFileAmplitudes [8302] = 8'd122;
   assign soundFileAmplitudes [8303] = 8'd131;
   assign soundFileAmplitudes [8304] = 8'd123;
   assign soundFileAmplitudes [8305] = 8'd127;
   assign soundFileAmplitudes [8306] = 8'd127;
   assign soundFileAmplitudes [8307] = 8'd121;
   assign soundFileAmplitudes [8308] = 8'd129;
   assign soundFileAmplitudes [8309] = 8'd110;
   assign soundFileAmplitudes [8310] = 8'd118;
   assign soundFileAmplitudes [8311] = 8'd142;
   assign soundFileAmplitudes [8312] = 8'd145;
   assign soundFileAmplitudes [8313] = 8'd144;
   assign soundFileAmplitudes [8314] = 8'd139;
   assign soundFileAmplitudes [8315] = 8'd136;
   assign soundFileAmplitudes [8316] = 8'd141;
   assign soundFileAmplitudes [8317] = 8'd140;
   assign soundFileAmplitudes [8318] = 8'd142;
   assign soundFileAmplitudes [8319] = 8'd143;
   assign soundFileAmplitudes [8320] = 8'd135;
   assign soundFileAmplitudes [8321] = 8'd120;
   assign soundFileAmplitudes [8322] = 8'd110;
   assign soundFileAmplitudes [8323] = 8'd112;
   assign soundFileAmplitudes [8324] = 8'd111;
   assign soundFileAmplitudes [8325] = 8'd116;
   assign soundFileAmplitudes [8326] = 8'd115;
   assign soundFileAmplitudes [8327] = 8'd107;
   assign soundFileAmplitudes [8328] = 8'd108;
   assign soundFileAmplitudes [8329] = 8'd124;
   assign soundFileAmplitudes [8330] = 8'd136;
   assign soundFileAmplitudes [8331] = 8'd148;
   assign soundFileAmplitudes [8332] = 8'd149;
   assign soundFileAmplitudes [8333] = 8'd139;
   assign soundFileAmplitudes [8334] = 8'd126;
   assign soundFileAmplitudes [8335] = 8'd115;
   assign soundFileAmplitudes [8336] = 8'd126;
   assign soundFileAmplitudes [8337] = 8'd118;
   assign soundFileAmplitudes [8338] = 8'd120;
   assign soundFileAmplitudes [8339] = 8'd115;
   assign soundFileAmplitudes [8340] = 8'd108;
   assign soundFileAmplitudes [8341] = 8'd114;
   assign soundFileAmplitudes [8342] = 8'd107;
   assign soundFileAmplitudes [8343] = 8'd113;
   assign soundFileAmplitudes [8344] = 8'd126;
   assign soundFileAmplitudes [8345] = 8'd127;
   assign soundFileAmplitudes [8346] = 8'd129;
   assign soundFileAmplitudes [8347] = 8'd142;
   assign soundFileAmplitudes [8348] = 8'd140;
   assign soundFileAmplitudes [8349] = 8'd143;
   assign soundFileAmplitudes [8350] = 8'd147;
   assign soundFileAmplitudes [8351] = 8'd150;
   assign soundFileAmplitudes [8352] = 8'd158;
   assign soundFileAmplitudes [8353] = 8'd139;
   assign soundFileAmplitudes [8354] = 8'd123;
   assign soundFileAmplitudes [8355] = 8'd118;
   assign soundFileAmplitudes [8356] = 8'd109;
   assign soundFileAmplitudes [8357] = 8'd114;
   assign soundFileAmplitudes [8358] = 8'd107;
   assign soundFileAmplitudes [8359] = 8'd95;
   assign soundFileAmplitudes [8360] = 8'd91;
   assign soundFileAmplitudes [8361] = 8'd95;
   assign soundFileAmplitudes [8362] = 8'd107;
   assign soundFileAmplitudes [8363] = 8'd116;
   assign soundFileAmplitudes [8364] = 8'd128;
   assign soundFileAmplitudes [8365] = 8'd141;
   assign soundFileAmplitudes [8366] = 8'd137;
   assign soundFileAmplitudes [8367] = 8'd135;
   assign soundFileAmplitudes [8368] = 8'd143;
   assign soundFileAmplitudes [8369] = 8'd146;
   assign soundFileAmplitudes [8370] = 8'd142;
   assign soundFileAmplitudes [8371] = 8'd136;
   assign soundFileAmplitudes [8372] = 8'd132;
   assign soundFileAmplitudes [8373] = 8'd125;
   assign soundFileAmplitudes [8374] = 8'd115;
   assign soundFileAmplitudes [8375] = 8'd113;
   assign soundFileAmplitudes [8376] = 8'd128;
   assign soundFileAmplitudes [8377] = 8'd132;
   assign soundFileAmplitudes [8378] = 8'd125;
   assign soundFileAmplitudes [8379] = 8'd122;
   assign soundFileAmplitudes [8380] = 8'd126;
   assign soundFileAmplitudes [8381] = 8'd129;
   assign soundFileAmplitudes [8382] = 8'd136;
   assign soundFileAmplitudes [8383] = 8'd148;
   assign soundFileAmplitudes [8384] = 8'd152;
   assign soundFileAmplitudes [8385] = 8'd148;
   assign soundFileAmplitudes [8386] = 8'd133;
   assign soundFileAmplitudes [8387] = 8'd127;
   assign soundFileAmplitudes [8388] = 8'd128;
   assign soundFileAmplitudes [8389] = 8'd130;
   assign soundFileAmplitudes [8390] = 8'd122;
   assign soundFileAmplitudes [8391] = 8'd108;
   assign soundFileAmplitudes [8392] = 8'd84;
   assign soundFileAmplitudes [8393] = 8'd78;
   assign soundFileAmplitudes [8394] = 8'd98;
   assign soundFileAmplitudes [8395] = 8'd111;
   assign soundFileAmplitudes [8396] = 8'd119;
   assign soundFileAmplitudes [8397] = 8'd117;
   assign soundFileAmplitudes [8398] = 8'd112;
   assign soundFileAmplitudes [8399] = 8'd101;
   assign soundFileAmplitudes [8400] = 8'd124;
   assign soundFileAmplitudes [8401] = 8'd145;
   assign soundFileAmplitudes [8402] = 8'd151;
   assign soundFileAmplitudes [8403] = 8'd160;
   assign soundFileAmplitudes [8404] = 8'd146;
   assign soundFileAmplitudes [8405] = 8'd150;
   assign soundFileAmplitudes [8406] = 8'd133;
   assign soundFileAmplitudes [8407] = 8'd124;
   assign soundFileAmplitudes [8408] = 8'd136;
   assign soundFileAmplitudes [8409] = 8'd146;
   assign soundFileAmplitudes [8410] = 8'd140;
   assign soundFileAmplitudes [8411] = 8'd127;
   assign soundFileAmplitudes [8412] = 8'd123;
   assign soundFileAmplitudes [8413] = 8'd122;
   assign soundFileAmplitudes [8414] = 8'd126;
   assign soundFileAmplitudes [8415] = 8'd126;
   assign soundFileAmplitudes [8416] = 8'd138;
   assign soundFileAmplitudes [8417] = 8'd144;
   assign soundFileAmplitudes [8418] = 8'd146;
   assign soundFileAmplitudes [8419] = 8'd134;
   assign soundFileAmplitudes [8420] = 8'd123;
   assign soundFileAmplitudes [8421] = 8'd119;
   assign soundFileAmplitudes [8422] = 8'd122;
   assign soundFileAmplitudes [8423] = 8'd123;
   assign soundFileAmplitudes [8424] = 8'd116;
   assign soundFileAmplitudes [8425] = 8'd107;
   assign soundFileAmplitudes [8426] = 8'd100;
   assign soundFileAmplitudes [8427] = 8'd101;
   assign soundFileAmplitudes [8428] = 8'd108;
   assign soundFileAmplitudes [8429] = 8'd120;
   assign soundFileAmplitudes [8430] = 8'd118;
   assign soundFileAmplitudes [8431] = 8'd119;
   assign soundFileAmplitudes [8432] = 8'd118;
   assign soundFileAmplitudes [8433] = 8'd126;
   assign soundFileAmplitudes [8434] = 8'd127;
   assign soundFileAmplitudes [8435] = 8'd129;
   assign soundFileAmplitudes [8436] = 8'd128;
   assign soundFileAmplitudes [8437] = 8'd130;
   assign soundFileAmplitudes [8438] = 8'd145;
   assign soundFileAmplitudes [8439] = 8'd133;
   assign soundFileAmplitudes [8440] = 8'd141;
   assign soundFileAmplitudes [8441] = 8'd150;
   assign soundFileAmplitudes [8442] = 8'd140;
   assign soundFileAmplitudes [8443] = 8'd128;
   assign soundFileAmplitudes [8444] = 8'd130;
   assign soundFileAmplitudes [8445] = 8'd134;
   assign soundFileAmplitudes [8446] = 8'd135;
   assign soundFileAmplitudes [8447] = 8'd140;
   assign soundFileAmplitudes [8448] = 8'd130;
   assign soundFileAmplitudes [8449] = 8'd140;
   assign soundFileAmplitudes [8450] = 8'd142;
   assign soundFileAmplitudes [8451] = 8'd127;
   assign soundFileAmplitudes [8452] = 8'd122;
   assign soundFileAmplitudes [8453] = 8'd124;
   assign soundFileAmplitudes [8454] = 8'd132;
   assign soundFileAmplitudes [8455] = 8'd140;
   assign soundFileAmplitudes [8456] = 8'd132;
   assign soundFileAmplitudes [8457] = 8'd121;
   assign soundFileAmplitudes [8458] = 8'd114;
   assign soundFileAmplitudes [8459] = 8'd109;
   assign soundFileAmplitudes [8460] = 8'd115;
   assign soundFileAmplitudes [8461] = 8'd126;
   assign soundFileAmplitudes [8462] = 8'd125;
   assign soundFileAmplitudes [8463] = 8'd111;
   assign soundFileAmplitudes [8464] = 8'd101;
   assign soundFileAmplitudes [8465] = 8'd111;
   assign soundFileAmplitudes [8466] = 8'd121;
   assign soundFileAmplitudes [8467] = 8'd121;
   assign soundFileAmplitudes [8468] = 8'd130;
   assign soundFileAmplitudes [8469] = 8'd121;
   assign soundFileAmplitudes [8470] = 8'd124;
   assign soundFileAmplitudes [8471] = 8'd114;
   assign soundFileAmplitudes [8472] = 8'd113;
   assign soundFileAmplitudes [8473] = 8'd135;
   assign soundFileAmplitudes [8474] = 8'd140;
   assign soundFileAmplitudes [8475] = 8'd140;
   assign soundFileAmplitudes [8476] = 8'd138;
   assign soundFileAmplitudes [8477] = 8'd140;
   assign soundFileAmplitudes [8478] = 8'd130;
   assign soundFileAmplitudes [8479] = 8'd123;
   assign soundFileAmplitudes [8480] = 8'd122;
   assign soundFileAmplitudes [8481] = 8'd125;
   assign soundFileAmplitudes [8482] = 8'd137;
   assign soundFileAmplitudes [8483] = 8'd140;
   assign soundFileAmplitudes [8484] = 8'd130;
   assign soundFileAmplitudes [8485] = 8'd122;
   assign soundFileAmplitudes [8486] = 8'd119;
   assign soundFileAmplitudes [8487] = 8'd123;
   assign soundFileAmplitudes [8488] = 8'd122;
   assign soundFileAmplitudes [8489] = 8'd121;
   assign soundFileAmplitudes [8490] = 8'd122;
   assign soundFileAmplitudes [8491] = 8'd129;
   assign soundFileAmplitudes [8492] = 8'd130;
   assign soundFileAmplitudes [8493] = 8'd130;
   assign soundFileAmplitudes [8494] = 8'd130;
   assign soundFileAmplitudes [8495] = 8'd124;
   assign soundFileAmplitudes [8496] = 8'd120;
   assign soundFileAmplitudes [8497] = 8'd123;
   assign soundFileAmplitudes [8498] = 8'd130;
   assign soundFileAmplitudes [8499] = 8'd118;
   assign soundFileAmplitudes [8500] = 8'd119;
   assign soundFileAmplitudes [8501] = 8'd117;
   assign soundFileAmplitudes [8502] = 8'd117;
   assign soundFileAmplitudes [8503] = 8'd126;
   assign soundFileAmplitudes [8504] = 8'd122;
   assign soundFileAmplitudes [8505] = 8'd126;
   assign soundFileAmplitudes [8506] = 8'd131;
   assign soundFileAmplitudes [8507] = 8'd125;
   assign soundFileAmplitudes [8508] = 8'd128;
   assign soundFileAmplitudes [8509] = 8'd135;
   assign soundFileAmplitudes [8510] = 8'd133;
   assign soundFileAmplitudes [8511] = 8'd132;
   assign soundFileAmplitudes [8512] = 8'd129;
   assign soundFileAmplitudes [8513] = 8'd133;
   assign soundFileAmplitudes [8514] = 8'd131;
   assign soundFileAmplitudes [8515] = 8'd131;
   assign soundFileAmplitudes [8516] = 8'd125;
   assign soundFileAmplitudes [8517] = 8'd113;
   assign soundFileAmplitudes [8518] = 8'd115;
   assign soundFileAmplitudes [8519] = 8'd119;
   assign soundFileAmplitudes [8520] = 8'd122;
   assign soundFileAmplitudes [8521] = 8'd126;
   assign soundFileAmplitudes [8522] = 8'd117;
   assign soundFileAmplitudes [8523] = 8'd112;
   assign soundFileAmplitudes [8524] = 8'd119;
   assign soundFileAmplitudes [8525] = 8'd122;
   assign soundFileAmplitudes [8526] = 8'd138;
   assign soundFileAmplitudes [8527] = 8'd142;
   assign soundFileAmplitudes [8528] = 8'd133;
   assign soundFileAmplitudes [8529] = 8'd121;
   assign soundFileAmplitudes [8530] = 8'd124;
   assign soundFileAmplitudes [8531] = 8'd134;
   assign soundFileAmplitudes [8532] = 8'd138;
   assign soundFileAmplitudes [8533] = 8'd141;
   assign soundFileAmplitudes [8534] = 8'd125;
   assign soundFileAmplitudes [8535] = 8'd117;
   assign soundFileAmplitudes [8536] = 8'd114;
   assign soundFileAmplitudes [8537] = 8'd117;
   assign soundFileAmplitudes [8538] = 8'd134;
   assign soundFileAmplitudes [8539] = 8'd142;
   assign soundFileAmplitudes [8540] = 8'd133;
   assign soundFileAmplitudes [8541] = 8'd126;
   assign soundFileAmplitudes [8542] = 8'd125;
   assign soundFileAmplitudes [8543] = 8'd125;
   assign soundFileAmplitudes [8544] = 8'd136;
   assign soundFileAmplitudes [8545] = 8'd143;
   assign soundFileAmplitudes [8546] = 8'd137;
   assign soundFileAmplitudes [8547] = 8'd129;
   assign soundFileAmplitudes [8548] = 8'd127;
   assign soundFileAmplitudes [8549] = 8'd121;
   assign soundFileAmplitudes [8550] = 8'd115;
   assign soundFileAmplitudes [8551] = 8'd121;
   assign soundFileAmplitudes [8552] = 8'd125;
   assign soundFileAmplitudes [8553] = 8'd124;
   assign soundFileAmplitudes [8554] = 8'd115;
   assign soundFileAmplitudes [8555] = 8'd109;
   assign soundFileAmplitudes [8556] = 8'd108;
   assign soundFileAmplitudes [8557] = 8'd115;
   assign soundFileAmplitudes [8558] = 8'd124;
   assign soundFileAmplitudes [8559] = 8'd129;
   assign soundFileAmplitudes [8560] = 8'd129;
   assign soundFileAmplitudes [8561] = 8'd126;
   assign soundFileAmplitudes [8562] = 8'd129;
   assign soundFileAmplitudes [8563] = 8'd132;
   assign soundFileAmplitudes [8564] = 8'd139;
   assign soundFileAmplitudes [8565] = 8'd139;
   assign soundFileAmplitudes [8566] = 8'd142;
   assign soundFileAmplitudes [8567] = 8'd136;
   assign soundFileAmplitudes [8568] = 8'd134;
   assign soundFileAmplitudes [8569] = 8'd133;
   assign soundFileAmplitudes [8570] = 8'd125;
   assign soundFileAmplitudes [8571] = 8'd126;
   assign soundFileAmplitudes [8572] = 8'd125;
   assign soundFileAmplitudes [8573] = 8'd125;
   assign soundFileAmplitudes [8574] = 8'd130;
   assign soundFileAmplitudes [8575] = 8'd134;
   assign soundFileAmplitudes [8576] = 8'd134;
   assign soundFileAmplitudes [8577] = 8'd135;
   assign soundFileAmplitudes [8578] = 8'd124;
   assign soundFileAmplitudes [8579] = 8'd129;
   assign soundFileAmplitudes [8580] = 8'd143;
   assign soundFileAmplitudes [8581] = 8'd142;
   assign soundFileAmplitudes [8582] = 8'd127;
   assign soundFileAmplitudes [8583] = 8'd120;
   assign soundFileAmplitudes [8584] = 8'd121;
   assign soundFileAmplitudes [8585] = 8'd107;
   assign soundFileAmplitudes [8586] = 8'd103;
   assign soundFileAmplitudes [8587] = 8'd106;
   assign soundFileAmplitudes [8588] = 8'd108;
   assign soundFileAmplitudes [8589] = 8'd112;
   assign soundFileAmplitudes [8590] = 8'd115;
   assign soundFileAmplitudes [8591] = 8'd117;
   assign soundFileAmplitudes [8592] = 8'd125;
   assign soundFileAmplitudes [8593] = 8'd120;
   assign soundFileAmplitudes [8594] = 8'd118;
   assign soundFileAmplitudes [8595] = 8'd122;
   assign soundFileAmplitudes [8596] = 8'd134;
   assign soundFileAmplitudes [8597] = 8'd149;
   assign soundFileAmplitudes [8598] = 8'd154;
   assign soundFileAmplitudes [8599] = 8'd154;
   assign soundFileAmplitudes [8600] = 8'd137;
   assign soundFileAmplitudes [8601] = 8'd135;
   assign soundFileAmplitudes [8602] = 8'd137;
   assign soundFileAmplitudes [8603] = 8'd136;
   assign soundFileAmplitudes [8604] = 8'd137;
   assign soundFileAmplitudes [8605] = 8'd127;
   assign soundFileAmplitudes [8606] = 8'd117;
   assign soundFileAmplitudes [8607] = 8'd109;
   assign soundFileAmplitudes [8608] = 8'd111;
   assign soundFileAmplitudes [8609] = 8'd121;
   assign soundFileAmplitudes [8610] = 8'd131;
   assign soundFileAmplitudes [8611] = 8'd130;
   assign soundFileAmplitudes [8612] = 8'd128;
   assign soundFileAmplitudes [8613] = 8'd119;
   assign soundFileAmplitudes [8614] = 8'd116;
   assign soundFileAmplitudes [8615] = 8'd127;
   assign soundFileAmplitudes [8616] = 8'd137;
   assign soundFileAmplitudes [8617] = 8'd140;
   assign soundFileAmplitudes [8618] = 8'd131;
   assign soundFileAmplitudes [8619] = 8'd126;
   assign soundFileAmplitudes [8620] = 8'd117;
   assign soundFileAmplitudes [8621] = 8'd107;
   assign soundFileAmplitudes [8622] = 8'd109;
   assign soundFileAmplitudes [8623] = 8'd111;
   assign soundFileAmplitudes [8624] = 8'd110;
   assign soundFileAmplitudes [8625] = 8'd117;
   assign soundFileAmplitudes [8626] = 8'd112;
   assign soundFileAmplitudes [8627] = 8'd115;
   assign soundFileAmplitudes [8628] = 8'd121;
   assign soundFileAmplitudes [8629] = 8'd121;
   assign soundFileAmplitudes [8630] = 8'd135;
   assign soundFileAmplitudes [8631] = 8'd135;
   assign soundFileAmplitudes [8632] = 8'd145;
   assign soundFileAmplitudes [8633] = 8'd153;
   assign soundFileAmplitudes [8634] = 8'd149;
   assign soundFileAmplitudes [8635] = 8'd148;
   assign soundFileAmplitudes [8636] = 8'd144;
   assign soundFileAmplitudes [8637] = 8'd137;
   assign soundFileAmplitudes [8638] = 8'd136;
   assign soundFileAmplitudes [8639] = 8'd130;
   assign soundFileAmplitudes [8640] = 8'd118;
   assign soundFileAmplitudes [8641] = 8'd117;
   assign soundFileAmplitudes [8642] = 8'd110;
   assign soundFileAmplitudes [8643] = 8'd109;
   assign soundFileAmplitudes [8644] = 8'd117;
   assign soundFileAmplitudes [8645] = 8'd116;
   assign soundFileAmplitudes [8646] = 8'd112;
   assign soundFileAmplitudes [8647] = 8'd115;
   assign soundFileAmplitudes [8648] = 8'd118;
   assign soundFileAmplitudes [8649] = 8'd123;
   assign soundFileAmplitudes [8650] = 8'd135;
   assign soundFileAmplitudes [8651] = 8'd139;
   assign soundFileAmplitudes [8652] = 8'd134;
   assign soundFileAmplitudes [8653] = 8'd125;
   assign soundFileAmplitudes [8654] = 8'd122;
   assign soundFileAmplitudes [8655] = 8'd115;
   assign soundFileAmplitudes [8656] = 8'd112;
   assign soundFileAmplitudes [8657] = 8'd116;
   assign soundFileAmplitudes [8658] = 8'd114;
   assign soundFileAmplitudes [8659] = 8'd112;
   assign soundFileAmplitudes [8660] = 8'd114;
   assign soundFileAmplitudes [8661] = 8'd109;
   assign soundFileAmplitudes [8662] = 8'd114;
   assign soundFileAmplitudes [8663] = 8'd132;
   assign soundFileAmplitudes [8664] = 8'd137;
   assign soundFileAmplitudes [8665] = 8'd139;
   assign soundFileAmplitudes [8666] = 8'd141;
   assign soundFileAmplitudes [8667] = 8'd147;
   assign soundFileAmplitudes [8668] = 8'd155;
   assign soundFileAmplitudes [8669] = 8'd165;
   assign soundFileAmplitudes [8670] = 8'd150;
   assign soundFileAmplitudes [8671] = 8'd139;
   assign soundFileAmplitudes [8672] = 8'd141;
   assign soundFileAmplitudes [8673] = 8'd135;
   assign soundFileAmplitudes [8674] = 8'd131;
   assign soundFileAmplitudes [8675] = 8'd120;
   assign soundFileAmplitudes [8676] = 8'd112;
   assign soundFileAmplitudes [8677] = 8'd105;
   assign soundFileAmplitudes [8678] = 8'd105;
   assign soundFileAmplitudes [8679] = 8'd106;
   assign soundFileAmplitudes [8680] = 8'd115;
   assign soundFileAmplitudes [8681] = 8'd122;
   assign soundFileAmplitudes [8682] = 8'd121;
   assign soundFileAmplitudes [8683] = 8'd113;
   assign soundFileAmplitudes [8684] = 8'd117;
   assign soundFileAmplitudes [8685] = 8'd133;
   assign soundFileAmplitudes [8686] = 8'd141;
   assign soundFileAmplitudes [8687] = 8'd137;
   assign soundFileAmplitudes [8688] = 8'd127;
   assign soundFileAmplitudes [8689] = 8'd131;
   assign soundFileAmplitudes [8690] = 8'd118;
   assign soundFileAmplitudes [8691] = 8'd114;
   assign soundFileAmplitudes [8692] = 8'd118;
   assign soundFileAmplitudes [8693] = 8'd116;
   assign soundFileAmplitudes [8694] = 8'd118;
   assign soundFileAmplitudes [8695] = 8'd120;
   assign soundFileAmplitudes [8696] = 8'd118;
   assign soundFileAmplitudes [8697] = 8'd113;
   assign soundFileAmplitudes [8698] = 8'd116;
   assign soundFileAmplitudes [8699] = 8'd125;
   assign soundFileAmplitudes [8700] = 8'd143;
   assign soundFileAmplitudes [8701] = 8'd151;
   assign soundFileAmplitudes [8702] = 8'd150;
   assign soundFileAmplitudes [8703] = 8'd154;
   assign soundFileAmplitudes [8704] = 8'd150;
   assign soundFileAmplitudes [8705] = 8'd144;
   assign soundFileAmplitudes [8706] = 8'd149;
   assign soundFileAmplitudes [8707] = 8'd149;
   assign soundFileAmplitudes [8708] = 8'd142;
   assign soundFileAmplitudes [8709] = 8'd134;
   assign soundFileAmplitudes [8710] = 8'd119;
   assign soundFileAmplitudes [8711] = 8'd102;
   assign soundFileAmplitudes [8712] = 8'd95;
   assign soundFileAmplitudes [8713] = 8'd97;
   assign soundFileAmplitudes [8714] = 8'd113;
   assign soundFileAmplitudes [8715] = 8'd126;
   assign soundFileAmplitudes [8716] = 8'd127;
   assign soundFileAmplitudes [8717] = 8'd118;
   assign soundFileAmplitudes [8718] = 8'd115;
   assign soundFileAmplitudes [8719] = 8'd132;
   assign soundFileAmplitudes [8720] = 8'd141;
   assign soundFileAmplitudes [8721] = 8'd146;
   assign soundFileAmplitudes [8722] = 8'd140;
   assign soundFileAmplitudes [8723] = 8'd133;
   assign soundFileAmplitudes [8724] = 8'd124;
   assign soundFileAmplitudes [8725] = 8'd109;
   assign soundFileAmplitudes [8726] = 8'd113;
   assign soundFileAmplitudes [8727] = 8'd124;
   assign soundFileAmplitudes [8728] = 8'd125;
   assign soundFileAmplitudes [8729] = 8'd117;
   assign soundFileAmplitudes [8730] = 8'd109;
   assign soundFileAmplitudes [8731] = 8'd110;
   assign soundFileAmplitudes [8732] = 8'd121;
   assign soundFileAmplitudes [8733] = 8'd124;
   assign soundFileAmplitudes [8734] = 8'd129;
   assign soundFileAmplitudes [8735] = 8'd130;
   assign soundFileAmplitudes [8736] = 8'd124;
   assign soundFileAmplitudes [8737] = 8'd141;
   assign soundFileAmplitudes [8738] = 8'd147;
   assign soundFileAmplitudes [8739] = 8'd142;
   assign soundFileAmplitudes [8740] = 8'd145;
   assign soundFileAmplitudes [8741] = 8'd145;
   assign soundFileAmplitudes [8742] = 8'd139;
   assign soundFileAmplitudes [8743] = 8'd131;
   assign soundFileAmplitudes [8744] = 8'd127;
   assign soundFileAmplitudes [8745] = 8'd113;
   assign soundFileAmplitudes [8746] = 8'd110;
   assign soundFileAmplitudes [8747] = 8'd108;
   assign soundFileAmplitudes [8748] = 8'd115;
   assign soundFileAmplitudes [8749] = 8'd128;
   assign soundFileAmplitudes [8750] = 8'd123;
   assign soundFileAmplitudes [8751] = 8'd119;
   assign soundFileAmplitudes [8752] = 8'd112;
   assign soundFileAmplitudes [8753] = 8'd134;
   assign soundFileAmplitudes [8754] = 8'd150;
   assign soundFileAmplitudes [8755] = 8'd149;
   assign soundFileAmplitudes [8756] = 8'd138;
   assign soundFileAmplitudes [8757] = 8'd125;
   assign soundFileAmplitudes [8758] = 8'd116;
   assign soundFileAmplitudes [8759] = 8'd108;
   assign soundFileAmplitudes [8760] = 8'd111;
   assign soundFileAmplitudes [8761] = 8'd117;
   assign soundFileAmplitudes [8762] = 8'd119;
   assign soundFileAmplitudes [8763] = 8'd119;
   assign soundFileAmplitudes [8764] = 8'd119;
   assign soundFileAmplitudes [8765] = 8'd118;
   assign soundFileAmplitudes [8766] = 8'd127;
   assign soundFileAmplitudes [8767] = 8'd132;
   assign soundFileAmplitudes [8768] = 8'd139;
   assign soundFileAmplitudes [8769] = 8'd140;
   assign soundFileAmplitudes [8770] = 8'd137;
   assign soundFileAmplitudes [8771] = 8'd132;
   assign soundFileAmplitudes [8772] = 8'd138;
   assign soundFileAmplitudes [8773] = 8'd139;
   assign soundFileAmplitudes [8774] = 8'd131;
   assign soundFileAmplitudes [8775] = 8'd133;
   assign soundFileAmplitudes [8776] = 8'd131;
   assign soundFileAmplitudes [8777] = 8'd125;
   assign soundFileAmplitudes [8778] = 8'd116;
   assign soundFileAmplitudes [8779] = 8'd105;
   assign soundFileAmplitudes [8780] = 8'd96;
   assign soundFileAmplitudes [8781] = 8'd99;
   assign soundFileAmplitudes [8782] = 8'd111;
   assign soundFileAmplitudes [8783] = 8'd123;
   assign soundFileAmplitudes [8784] = 8'd125;
   assign soundFileAmplitudes [8785] = 8'd124;
   assign soundFileAmplitudes [8786] = 8'd120;
   assign soundFileAmplitudes [8787] = 8'd118;
   assign soundFileAmplitudes [8788] = 8'd136;
   assign soundFileAmplitudes [8789] = 8'd148;
   assign soundFileAmplitudes [8790] = 8'd139;
   assign soundFileAmplitudes [8791] = 8'd132;
   assign soundFileAmplitudes [8792] = 8'd130;
   assign soundFileAmplitudes [8793] = 8'd114;
   assign soundFileAmplitudes [8794] = 8'd110;
   assign soundFileAmplitudes [8795] = 8'd119;
   assign soundFileAmplitudes [8796] = 8'd126;
   assign soundFileAmplitudes [8797] = 8'd129;
   assign soundFileAmplitudes [8798] = 8'd134;
   assign soundFileAmplitudes [8799] = 8'd130;
   assign soundFileAmplitudes [8800] = 8'd128;
   assign soundFileAmplitudes [8801] = 8'd137;
   assign soundFileAmplitudes [8802] = 8'd137;
   assign soundFileAmplitudes [8803] = 8'd143;
   assign soundFileAmplitudes [8804] = 8'd141;
   assign soundFileAmplitudes [8805] = 8'd137;
   assign soundFileAmplitudes [8806] = 8'd135;
   assign soundFileAmplitudes [8807] = 8'd143;
   assign soundFileAmplitudes [8808] = 8'd131;
   assign soundFileAmplitudes [8809] = 8'd114;
   assign soundFileAmplitudes [8810] = 8'd117;
   assign soundFileAmplitudes [8811] = 8'd120;
   assign soundFileAmplitudes [8812] = 8'd123;
   assign soundFileAmplitudes [8813] = 8'd114;
   assign soundFileAmplitudes [8814] = 8'd107;
   assign soundFileAmplitudes [8815] = 8'd101;
   assign soundFileAmplitudes [8816] = 8'd107;
   assign soundFileAmplitudes [8817] = 8'd125;
   assign soundFileAmplitudes [8818] = 8'd133;
   assign soundFileAmplitudes [8819] = 8'd132;
   assign soundFileAmplitudes [8820] = 8'd128;
   assign soundFileAmplitudes [8821] = 8'd119;
   assign soundFileAmplitudes [8822] = 8'd132;
   assign soundFileAmplitudes [8823] = 8'd148;
   assign soundFileAmplitudes [8824] = 8'd142;
   assign soundFileAmplitudes [8825] = 8'd125;
   assign soundFileAmplitudes [8826] = 8'd120;
   assign soundFileAmplitudes [8827] = 8'd119;
   assign soundFileAmplitudes [8828] = 8'd108;
   assign soundFileAmplitudes [8829] = 8'd114;
   assign soundFileAmplitudes [8830] = 8'd120;
   assign soundFileAmplitudes [8831] = 8'd121;
   assign soundFileAmplitudes [8832] = 8'd131;
   assign soundFileAmplitudes [8833] = 8'd134;
   assign soundFileAmplitudes [8834] = 8'd129;
   assign soundFileAmplitudes [8835] = 8'd138;
   assign soundFileAmplitudes [8836] = 8'd137;
   assign soundFileAmplitudes [8837] = 8'd141;
   assign soundFileAmplitudes [8838] = 8'd143;
   assign soundFileAmplitudes [8839] = 8'd139;
   assign soundFileAmplitudes [8840] = 8'd145;
   assign soundFileAmplitudes [8841] = 8'd137;
   assign soundFileAmplitudes [8842] = 8'd141;
   assign soundFileAmplitudes [8843] = 8'd133;
   assign soundFileAmplitudes [8844] = 8'd124;
   assign soundFileAmplitudes [8845] = 8'd126;
   assign soundFileAmplitudes [8846] = 8'd122;
   assign soundFileAmplitudes [8847] = 8'd116;
   assign soundFileAmplitudes [8848] = 8'd111;
   assign soundFileAmplitudes [8849] = 8'd106;
   assign soundFileAmplitudes [8850] = 8'd108;
   assign soundFileAmplitudes [8851] = 8'd129;
   assign soundFileAmplitudes [8852] = 8'd126;
   assign soundFileAmplitudes [8853] = 8'd122;
   assign soundFileAmplitudes [8854] = 8'd120;
   assign soundFileAmplitudes [8855] = 8'd120;
   assign soundFileAmplitudes [8856] = 8'd139;
   assign soundFileAmplitudes [8857] = 8'd153;
   assign soundFileAmplitudes [8858] = 8'd155;
   assign soundFileAmplitudes [8859] = 8'd141;
   assign soundFileAmplitudes [8860] = 8'd125;
   assign soundFileAmplitudes [8861] = 8'd112;
   assign soundFileAmplitudes [8862] = 8'd103;
   assign soundFileAmplitudes [8863] = 8'd105;
   assign soundFileAmplitudes [8864] = 8'd112;
   assign soundFileAmplitudes [8865] = 8'd113;
   assign soundFileAmplitudes [8866] = 8'd124;
   assign soundFileAmplitudes [8867] = 8'd123;
   assign soundFileAmplitudes [8868] = 8'd114;
   assign soundFileAmplitudes [8869] = 8'd118;
   assign soundFileAmplitudes [8870] = 8'd117;
   assign soundFileAmplitudes [8871] = 8'd125;
   assign soundFileAmplitudes [8872] = 8'd140;
   assign soundFileAmplitudes [8873] = 8'd149;
   assign soundFileAmplitudes [8874] = 8'd154;
   assign soundFileAmplitudes [8875] = 8'd148;
   assign soundFileAmplitudes [8876] = 8'd143;
   assign soundFileAmplitudes [8877] = 8'd146;
   assign soundFileAmplitudes [8878] = 8'd137;
   assign soundFileAmplitudes [8879] = 8'd127;
   assign soundFileAmplitudes [8880] = 8'd126;
   assign soundFileAmplitudes [8881] = 8'd124;
   assign soundFileAmplitudes [8882] = 8'd116;
   assign soundFileAmplitudes [8883] = 8'd93;
   assign soundFileAmplitudes [8884] = 8'd74;
   assign soundFileAmplitudes [8885] = 8'd93;
   assign soundFileAmplitudes [8886] = 8'd115;
   assign soundFileAmplitudes [8887] = 8'd125;
   assign soundFileAmplitudes [8888] = 8'd130;
   assign soundFileAmplitudes [8889] = 8'd129;
   assign soundFileAmplitudes [8890] = 8'd132;
   assign soundFileAmplitudes [8891] = 8'd147;
   assign soundFileAmplitudes [8892] = 8'd162;
   assign soundFileAmplitudes [8893] = 8'd149;
   assign soundFileAmplitudes [8894] = 8'd134;
   assign soundFileAmplitudes [8895] = 8'd135;
   assign soundFileAmplitudes [8896] = 8'd123;
   assign soundFileAmplitudes [8897] = 8'd110;
   assign soundFileAmplitudes [8898] = 8'd105;
   assign soundFileAmplitudes [8899] = 8'd102;
   assign soundFileAmplitudes [8900] = 8'd106;
   assign soundFileAmplitudes [8901] = 8'd114;
   assign soundFileAmplitudes [8902] = 8'd121;
   assign soundFileAmplitudes [8903] = 8'd126;
   assign soundFileAmplitudes [8904] = 8'd130;
   assign soundFileAmplitudes [8905] = 8'd128;
   assign soundFileAmplitudes [8906] = 8'd133;
   assign soundFileAmplitudes [8907] = 8'd144;
   assign soundFileAmplitudes [8908] = 8'd161;
   assign soundFileAmplitudes [8909] = 8'd158;
   assign soundFileAmplitudes [8910] = 8'd140;
   assign soundFileAmplitudes [8911] = 8'd145;
   assign soundFileAmplitudes [8912] = 8'd141;
   assign soundFileAmplitudes [8913] = 8'd124;
   assign soundFileAmplitudes [8914] = 8'd114;
   assign soundFileAmplitudes [8915] = 8'd108;
   assign soundFileAmplitudes [8916] = 8'd104;
   assign soundFileAmplitudes [8917] = 8'd95;
   assign soundFileAmplitudes [8918] = 8'd89;
   assign soundFileAmplitudes [8919] = 8'd94;
   assign soundFileAmplitudes [8920] = 8'd112;
   assign soundFileAmplitudes [8921] = 8'd130;
   assign soundFileAmplitudes [8922] = 8'd136;
   assign soundFileAmplitudes [8923] = 8'd135;
   assign soundFileAmplitudes [8924] = 8'd128;
   assign soundFileAmplitudes [8925] = 8'd142;
   assign soundFileAmplitudes [8926] = 8'd156;
   assign soundFileAmplitudes [8927] = 8'd151;
   assign soundFileAmplitudes [8928] = 8'd137;
   assign soundFileAmplitudes [8929] = 8'd127;
   assign soundFileAmplitudes [8930] = 8'd122;
   assign soundFileAmplitudes [8931] = 8'd100;
   assign soundFileAmplitudes [8932] = 8'd111;
   assign soundFileAmplitudes [8933] = 8'd119;
   assign soundFileAmplitudes [8934] = 8'd130;
   assign soundFileAmplitudes [8935] = 8'd134;
   assign soundFileAmplitudes [8936] = 8'd122;
   assign soundFileAmplitudes [8937] = 8'd122;
   assign soundFileAmplitudes [8938] = 8'd127;
   assign soundFileAmplitudes [8939] = 8'd127;
   assign soundFileAmplitudes [8940] = 8'd134;
   assign soundFileAmplitudes [8941] = 8'd140;
   assign soundFileAmplitudes [8942] = 8'd144;
   assign soundFileAmplitudes [8943] = 8'd147;
   assign soundFileAmplitudes [8944] = 8'd113;
   assign soundFileAmplitudes [8945] = 8'd123;
   assign soundFileAmplitudes [8946] = 8'd131;
   assign soundFileAmplitudes [8947] = 8'd122;
   assign soundFileAmplitudes [8948] = 8'd130;
   assign soundFileAmplitudes [8949] = 8'd124;
   assign soundFileAmplitudes [8950] = 8'd118;
   assign soundFileAmplitudes [8951] = 8'd117;
   assign soundFileAmplitudes [8952] = 8'd112;
   assign soundFileAmplitudes [8953] = 8'd103;
   assign soundFileAmplitudes [8954] = 8'd112;
   assign soundFileAmplitudes [8955] = 8'd130;
   assign soundFileAmplitudes [8956] = 8'd134;
   assign soundFileAmplitudes [8957] = 8'd131;
   assign soundFileAmplitudes [8958] = 8'd113;
   assign soundFileAmplitudes [8959] = 8'd117;
   assign soundFileAmplitudes [8960] = 8'd128;
   assign soundFileAmplitudes [8961] = 8'd126;
   assign soundFileAmplitudes [8962] = 8'd141;
   assign soundFileAmplitudes [8963] = 8'd136;
   assign soundFileAmplitudes [8964] = 8'd148;
   assign soundFileAmplitudes [8965] = 8'd129;
   assign soundFileAmplitudes [8966] = 8'd109;
   assign soundFileAmplitudes [8967] = 8'd127;
   assign soundFileAmplitudes [8968] = 8'd140;
   assign soundFileAmplitudes [8969] = 8'd146;
   assign soundFileAmplitudes [8970] = 8'd137;
   assign soundFileAmplitudes [8971] = 8'd135;
   assign soundFileAmplitudes [8972] = 8'd136;
   assign soundFileAmplitudes [8973] = 8'd128;
   assign soundFileAmplitudes [8974] = 8'd114;
   assign soundFileAmplitudes [8975] = 8'd124;
   assign soundFileAmplitudes [8976] = 8'd134;
   assign soundFileAmplitudes [8977] = 8'd134;
   assign soundFileAmplitudes [8978] = 8'd124;
   assign soundFileAmplitudes [8979] = 8'd123;
   assign soundFileAmplitudes [8980] = 8'd118;
   assign soundFileAmplitudes [8981] = 8'd124;
   assign soundFileAmplitudes [8982] = 8'd134;
   assign soundFileAmplitudes [8983] = 8'd131;
   assign soundFileAmplitudes [8984] = 8'd126;
   assign soundFileAmplitudes [8985] = 8'd118;
   assign soundFileAmplitudes [8986] = 8'd111;
   assign soundFileAmplitudes [8987] = 8'd104;
   assign soundFileAmplitudes [8988] = 8'd109;
   assign soundFileAmplitudes [8989] = 8'd116;
   assign soundFileAmplitudes [8990] = 8'd128;
   assign soundFileAmplitudes [8991] = 8'd125;
   assign soundFileAmplitudes [8992] = 8'd125;
   assign soundFileAmplitudes [8993] = 8'd120;
   assign soundFileAmplitudes [8994] = 8'd132;
   assign soundFileAmplitudes [8995] = 8'd144;
   assign soundFileAmplitudes [8996] = 8'd143;
   assign soundFileAmplitudes [8997] = 8'd145;
   assign soundFileAmplitudes [8998] = 8'd142;
   assign soundFileAmplitudes [8999] = 8'd142;
   assign soundFileAmplitudes [9000] = 8'd124;
   assign soundFileAmplitudes [9001] = 8'd122;
   assign soundFileAmplitudes [9002] = 8'd137;
   assign soundFileAmplitudes [9003] = 8'd143;
   assign soundFileAmplitudes [9004] = 8'd132;
   assign soundFileAmplitudes [9005] = 8'd115;
   assign soundFileAmplitudes [9006] = 8'd119;
   assign soundFileAmplitudes [9007] = 8'd127;
   assign soundFileAmplitudes [9008] = 8'd128;
   assign soundFileAmplitudes [9009] = 8'd118;
   assign soundFileAmplitudes [9010] = 8'd115;
   assign soundFileAmplitudes [9011] = 8'd126;
   assign soundFileAmplitudes [9012] = 8'd134;
   assign soundFileAmplitudes [9013] = 8'd143;
   assign soundFileAmplitudes [9014] = 8'd121;
   assign soundFileAmplitudes [9015] = 8'd108;
   assign soundFileAmplitudes [9016] = 8'd113;
   assign soundFileAmplitudes [9017] = 8'd121;
   assign soundFileAmplitudes [9018] = 8'd127;
   assign soundFileAmplitudes [9019] = 8'd110;
   assign soundFileAmplitudes [9020] = 8'd102;
   assign soundFileAmplitudes [9021] = 8'd94;
   assign soundFileAmplitudes [9022] = 8'd91;
   assign soundFileAmplitudes [9023] = 8'd113;
   assign soundFileAmplitudes [9024] = 8'd138;
   assign soundFileAmplitudes [9025] = 8'd151;
   assign soundFileAmplitudes [9026] = 8'd149;
   assign soundFileAmplitudes [9027] = 8'd139;
   assign soundFileAmplitudes [9028] = 8'd138;
   assign soundFileAmplitudes [9029] = 8'd152;
   assign soundFileAmplitudes [9030] = 8'd151;
   assign soundFileAmplitudes [9031] = 8'd137;
   assign soundFileAmplitudes [9032] = 8'd129;
   assign soundFileAmplitudes [9033] = 8'd128;
   assign soundFileAmplitudes [9034] = 8'd127;
   assign soundFileAmplitudes [9035] = 8'd101;
   assign soundFileAmplitudes [9036] = 8'd106;
   assign soundFileAmplitudes [9037] = 8'd123;
   assign soundFileAmplitudes [9038] = 8'd123;
   assign soundFileAmplitudes [9039] = 8'd119;
   assign soundFileAmplitudes [9040] = 8'd106;
   assign soundFileAmplitudes [9041] = 8'd117;
   assign soundFileAmplitudes [9042] = 8'd142;
   assign soundFileAmplitudes [9043] = 8'd146;
   assign soundFileAmplitudes [9044] = 8'd138;
   assign soundFileAmplitudes [9045] = 8'd125;
   assign soundFileAmplitudes [9046] = 8'd117;
   assign soundFileAmplitudes [9047] = 8'd129;
   assign soundFileAmplitudes [9048] = 8'd126;
   assign soundFileAmplitudes [9049] = 8'd123;
   assign soundFileAmplitudes [9050] = 8'd119;
   assign soundFileAmplitudes [9051] = 8'd118;
   assign soundFileAmplitudes [9052] = 8'd108;
   assign soundFileAmplitudes [9053] = 8'd101;
   assign soundFileAmplitudes [9054] = 8'd117;
   assign soundFileAmplitudes [9055] = 8'd122;
   assign soundFileAmplitudes [9056] = 8'd124;
   assign soundFileAmplitudes [9057] = 8'd117;
   assign soundFileAmplitudes [9058] = 8'd120;
   assign soundFileAmplitudes [9059] = 8'd137;
   assign soundFileAmplitudes [9060] = 8'd159;
   assign soundFileAmplitudes [9061] = 8'd157;
   assign soundFileAmplitudes [9062] = 8'd144;
   assign soundFileAmplitudes [9063] = 8'd138;
   assign soundFileAmplitudes [9064] = 8'd143;
   assign soundFileAmplitudes [9065] = 8'd143;
   assign soundFileAmplitudes [9066] = 8'd120;
   assign soundFileAmplitudes [9067] = 8'd118;
   assign soundFileAmplitudes [9068] = 8'd117;
   assign soundFileAmplitudes [9069] = 8'd108;
   assign soundFileAmplitudes [9070] = 8'd92;
   assign soundFileAmplitudes [9071] = 8'd98;
   assign soundFileAmplitudes [9072] = 8'd121;
   assign soundFileAmplitudes [9073] = 8'd129;
   assign soundFileAmplitudes [9074] = 8'd134;
   assign soundFileAmplitudes [9075] = 8'd136;
   assign soundFileAmplitudes [9076] = 8'd138;
   assign soundFileAmplitudes [9077] = 8'd138;
   assign soundFileAmplitudes [9078] = 8'd144;
   assign soundFileAmplitudes [9079] = 8'd138;
   assign soundFileAmplitudes [9080] = 8'd133;
   assign soundFileAmplitudes [9081] = 8'd138;
   assign soundFileAmplitudes [9082] = 8'd124;
   assign soundFileAmplitudes [9083] = 8'd112;
   assign soundFileAmplitudes [9084] = 8'd109;
   assign soundFileAmplitudes [9085] = 8'd119;
   assign soundFileAmplitudes [9086] = 8'd126;
   assign soundFileAmplitudes [9087] = 8'd125;
   assign soundFileAmplitudes [9088] = 8'd122;
   assign soundFileAmplitudes [9089] = 8'd121;
   assign soundFileAmplitudes [9090] = 8'd123;
   assign soundFileAmplitudes [9091] = 8'd130;
   assign soundFileAmplitudes [9092] = 8'd120;
   assign soundFileAmplitudes [9093] = 8'd126;
   assign soundFileAmplitudes [9094] = 8'd145;
   assign soundFileAmplitudes [9095] = 8'd149;
   assign soundFileAmplitudes [9096] = 8'd139;
   assign soundFileAmplitudes [9097] = 8'd113;
   assign soundFileAmplitudes [9098] = 8'd118;
   assign soundFileAmplitudes [9099] = 8'd133;
   assign soundFileAmplitudes [9100] = 8'd138;
   assign soundFileAmplitudes [9101] = 8'd131;
   assign soundFileAmplitudes [9102] = 8'd116;
   assign soundFileAmplitudes [9103] = 8'd116;
   assign soundFileAmplitudes [9104] = 8'd125;
   assign soundFileAmplitudes [9105] = 8'd126;
   assign soundFileAmplitudes [9106] = 8'd125;
   assign soundFileAmplitudes [9107] = 8'd117;
   assign soundFileAmplitudes [9108] = 8'd115;
   assign soundFileAmplitudes [9109] = 8'd132;
   assign soundFileAmplitudes [9110] = 8'd137;
   assign soundFileAmplitudes [9111] = 8'd126;
   assign soundFileAmplitudes [9112] = 8'd126;
   assign soundFileAmplitudes [9113] = 8'd117;
   assign soundFileAmplitudes [9114] = 8'd107;
   assign soundFileAmplitudes [9115] = 8'd122;
   assign soundFileAmplitudes [9116] = 8'd133;
   assign soundFileAmplitudes [9117] = 8'd142;
   assign soundFileAmplitudes [9118] = 8'd149;
   assign soundFileAmplitudes [9119] = 8'd136;
   assign soundFileAmplitudes [9120] = 8'd127;
   assign soundFileAmplitudes [9121] = 8'd129;
   assign soundFileAmplitudes [9122] = 8'd147;
   assign soundFileAmplitudes [9123] = 8'd139;
   assign soundFileAmplitudes [9124] = 8'd135;
   assign soundFileAmplitudes [9125] = 8'd129;
   assign soundFileAmplitudes [9126] = 8'd126;
   assign soundFileAmplitudes [9127] = 8'd119;
   assign soundFileAmplitudes [9128] = 8'd90;
   assign soundFileAmplitudes [9129] = 8'd107;
   assign soundFileAmplitudes [9130] = 8'd119;
   assign soundFileAmplitudes [9131] = 8'd121;
   assign soundFileAmplitudes [9132] = 8'd115;
   assign soundFileAmplitudes [9133] = 8'd111;
   assign soundFileAmplitudes [9134] = 8'd128;
   assign soundFileAmplitudes [9135] = 8'd144;
   assign soundFileAmplitudes [9136] = 8'd152;
   assign soundFileAmplitudes [9137] = 8'd143;
   assign soundFileAmplitudes [9138] = 8'd131;
   assign soundFileAmplitudes [9139] = 8'd138;
   assign soundFileAmplitudes [9140] = 8'd127;
   assign soundFileAmplitudes [9141] = 8'd118;
   assign soundFileAmplitudes [9142] = 8'd121;
   assign soundFileAmplitudes [9143] = 8'd120;
   assign soundFileAmplitudes [9144] = 8'd119;
   assign soundFileAmplitudes [9145] = 8'd97;
   assign soundFileAmplitudes [9146] = 8'd102;
   assign soundFileAmplitudes [9147] = 8'd117;
   assign soundFileAmplitudes [9148] = 8'd126;
   assign soundFileAmplitudes [9149] = 8'd132;
   assign soundFileAmplitudes [9150] = 8'd123;
   assign soundFileAmplitudes [9151] = 8'd128;
   assign soundFileAmplitudes [9152] = 8'd138;
   assign soundFileAmplitudes [9153] = 8'd153;
   assign soundFileAmplitudes [9154] = 8'd150;
   assign soundFileAmplitudes [9155] = 8'd141;
   assign soundFileAmplitudes [9156] = 8'd137;
   assign soundFileAmplitudes [9157] = 8'd140;
   assign soundFileAmplitudes [9158] = 8'd142;
   assign soundFileAmplitudes [9159] = 8'd114;
   assign soundFileAmplitudes [9160] = 8'd104;
   assign soundFileAmplitudes [9161] = 8'd101;
   assign soundFileAmplitudes [9162] = 8'd106;
   assign soundFileAmplitudes [9163] = 8'd113;
   assign soundFileAmplitudes [9164] = 8'd117;
   assign soundFileAmplitudes [9165] = 8'd119;
   assign soundFileAmplitudes [9166] = 8'd123;
   assign soundFileAmplitudes [9167] = 8'd131;
   assign soundFileAmplitudes [9168] = 8'd128;
   assign soundFileAmplitudes [9169] = 8'd134;
   assign soundFileAmplitudes [9170] = 8'd149;
   assign soundFileAmplitudes [9171] = 8'd148;
   assign soundFileAmplitudes [9172] = 8'd144;
   assign soundFileAmplitudes [9173] = 8'd139;
   assign soundFileAmplitudes [9174] = 8'd130;
   assign soundFileAmplitudes [9175] = 8'd115;
   assign soundFileAmplitudes [9176] = 8'd93;
   assign soundFileAmplitudes [9177] = 8'd106;
   assign soundFileAmplitudes [9178] = 8'd122;
   assign soundFileAmplitudes [9179] = 8'd124;
   assign soundFileAmplitudes [9180] = 8'd118;
   assign soundFileAmplitudes [9181] = 8'd107;
   assign soundFileAmplitudes [9182] = 8'd105;
   assign soundFileAmplitudes [9183] = 8'd108;
   assign soundFileAmplitudes [9184] = 8'd111;
   assign soundFileAmplitudes [9185] = 8'd129;
   assign soundFileAmplitudes [9186] = 8'd141;
   assign soundFileAmplitudes [9187] = 8'd145;
   assign soundFileAmplitudes [9188] = 8'd147;
   assign soundFileAmplitudes [9189] = 8'd136;
   assign soundFileAmplitudes [9190] = 8'd123;
   assign soundFileAmplitudes [9191] = 8'd121;
   assign soundFileAmplitudes [9192] = 8'd138;
   assign soundFileAmplitudes [9193] = 8'd143;
   assign soundFileAmplitudes [9194] = 8'd135;
   assign soundFileAmplitudes [9195] = 8'd119;
   assign soundFileAmplitudes [9196] = 8'd117;
   assign soundFileAmplitudes [9197] = 8'd128;
   assign soundFileAmplitudes [9198] = 8'd133;
   assign soundFileAmplitudes [9199] = 8'd131;
   assign soundFileAmplitudes [9200] = 8'd125;
   assign soundFileAmplitudes [9201] = 8'd131;
   assign soundFileAmplitudes [9202] = 8'd125;
   assign soundFileAmplitudes [9203] = 8'd119;
   assign soundFileAmplitudes [9204] = 8'd126;
   assign soundFileAmplitudes [9205] = 8'd129;
   assign soundFileAmplitudes [9206] = 8'd133;
   assign soundFileAmplitudes [9207] = 8'd129;
   assign soundFileAmplitudes [9208] = 8'd130;
   assign soundFileAmplitudes [9209] = 8'd134;
   assign soundFileAmplitudes [9210] = 8'd122;
   assign soundFileAmplitudes [9211] = 8'd120;
   assign soundFileAmplitudes [9212] = 8'd130;
   assign soundFileAmplitudes [9213] = 8'd122;
   assign soundFileAmplitudes [9214] = 8'd117;
   assign soundFileAmplitudes [9215] = 8'd119;
   assign soundFileAmplitudes [9216] = 8'd110;
   assign soundFileAmplitudes [9217] = 8'd123;
   assign soundFileAmplitudes [9218] = 8'd115;
   assign soundFileAmplitudes [9219] = 8'd101;
   assign soundFileAmplitudes [9220] = 8'd102;
   assign soundFileAmplitudes [9221] = 8'd106;
   assign soundFileAmplitudes [9222] = 8'd124;
   assign soundFileAmplitudes [9223] = 8'd137;
   assign soundFileAmplitudes [9224] = 8'd139;
   assign soundFileAmplitudes [9225] = 8'd131;
   assign soundFileAmplitudes [9226] = 8'd139;
   assign soundFileAmplitudes [9227] = 8'd143;
   assign soundFileAmplitudes [9228] = 8'd148;
   assign soundFileAmplitudes [9229] = 8'd153;
   assign soundFileAmplitudes [9230] = 8'd140;
   assign soundFileAmplitudes [9231] = 8'd124;
   assign soundFileAmplitudes [9232] = 8'd126;
   assign soundFileAmplitudes [9233] = 8'd130;
   assign soundFileAmplitudes [9234] = 8'd126;
   assign soundFileAmplitudes [9235] = 8'd123;
   assign soundFileAmplitudes [9236] = 8'd120;
   assign soundFileAmplitudes [9237] = 8'd120;
   assign soundFileAmplitudes [9238] = 8'd108;
   assign soundFileAmplitudes [9239] = 8'd114;
   assign soundFileAmplitudes [9240] = 8'd129;
   assign soundFileAmplitudes [9241] = 8'd142;
   assign soundFileAmplitudes [9242] = 8'd154;
   assign soundFileAmplitudes [9243] = 8'd146;
   assign soundFileAmplitudes [9244] = 8'd139;
   assign soundFileAmplitudes [9245] = 8'd130;
   assign soundFileAmplitudes [9246] = 8'd128;
   assign soundFileAmplitudes [9247] = 8'd135;
   assign soundFileAmplitudes [9248] = 8'd136;
   assign soundFileAmplitudes [9249] = 8'd126;
   assign soundFileAmplitudes [9250] = 8'd110;
   assign soundFileAmplitudes [9251] = 8'd93;
   assign soundFileAmplitudes [9252] = 8'd98;
   assign soundFileAmplitudes [9253] = 8'd97;
   assign soundFileAmplitudes [9254] = 8'd100;
   assign soundFileAmplitudes [9255] = 8'd110;
   assign soundFileAmplitudes [9256] = 8'd108;
   assign soundFileAmplitudes [9257] = 8'd126;
   assign soundFileAmplitudes [9258] = 8'd130;
   assign soundFileAmplitudes [9259] = 8'd133;
   assign soundFileAmplitudes [9260] = 8'd150;
   assign soundFileAmplitudes [9261] = 8'd149;
   assign soundFileAmplitudes [9262] = 8'd145;
   assign soundFileAmplitudes [9263] = 8'd154;
   assign soundFileAmplitudes [9264] = 8'd155;
   assign soundFileAmplitudes [9265] = 8'd147;
   assign soundFileAmplitudes [9266] = 8'd129;
   assign soundFileAmplitudes [9267] = 8'd119;
   assign soundFileAmplitudes [9268] = 8'd112;
   assign soundFileAmplitudes [9269] = 8'd110;
   assign soundFileAmplitudes [9270] = 8'd128;
   assign soundFileAmplitudes [9271] = 8'd140;
   assign soundFileAmplitudes [9272] = 8'd134;
   assign soundFileAmplitudes [9273] = 8'd123;
   assign soundFileAmplitudes [9274] = 8'd113;
   assign soundFileAmplitudes [9275] = 8'd127;
   assign soundFileAmplitudes [9276] = 8'd148;
   assign soundFileAmplitudes [9277] = 8'd149;
   assign soundFileAmplitudes [9278] = 8'd149;
   assign soundFileAmplitudes [9279] = 8'd138;
   assign soundFileAmplitudes [9280] = 8'd114;
   assign soundFileAmplitudes [9281] = 8'd90;
   assign soundFileAmplitudes [9282] = 8'd99;
   assign soundFileAmplitudes [9283] = 8'd107;
   assign soundFileAmplitudes [9284] = 8'd112;
   assign soundFileAmplitudes [9285] = 8'd106;
   assign soundFileAmplitudes [9286] = 8'd102;
   assign soundFileAmplitudes [9287] = 8'd105;
   assign soundFileAmplitudes [9288] = 8'd105;
   assign soundFileAmplitudes [9289] = 8'd124;
   assign soundFileAmplitudes [9290] = 8'd129;
   assign soundFileAmplitudes [9291] = 8'd119;
   assign soundFileAmplitudes [9292] = 8'd132;
   assign soundFileAmplitudes [9293] = 8'd146;
   assign soundFileAmplitudes [9294] = 8'd145;
   assign soundFileAmplitudes [9295] = 8'd141;
   assign soundFileAmplitudes [9296] = 8'd131;
   assign soundFileAmplitudes [9297] = 8'd129;
   assign soundFileAmplitudes [9298] = 8'd127;
   assign soundFileAmplitudes [9299] = 8'd126;
   assign soundFileAmplitudes [9300] = 8'd134;
   assign soundFileAmplitudes [9301] = 8'd137;
   assign soundFileAmplitudes [9302] = 8'd129;
   assign soundFileAmplitudes [9303] = 8'd132;
   assign soundFileAmplitudes [9304] = 8'd137;
   assign soundFileAmplitudes [9305] = 8'd150;
   assign soundFileAmplitudes [9306] = 8'd145;
   assign soundFileAmplitudes [9307] = 8'd136;
   assign soundFileAmplitudes [9308] = 8'd138;
   assign soundFileAmplitudes [9309] = 8'd133;
   assign soundFileAmplitudes [9310] = 8'd123;
   assign soundFileAmplitudes [9311] = 8'd111;
   assign soundFileAmplitudes [9312] = 8'd120;
   assign soundFileAmplitudes [9313] = 8'd114;
   assign soundFileAmplitudes [9314] = 8'd107;
   assign soundFileAmplitudes [9315] = 8'd101;
   assign soundFileAmplitudes [9316] = 8'd88;
   assign soundFileAmplitudes [9317] = 8'd97;
   assign soundFileAmplitudes [9318] = 8'd117;
   assign soundFileAmplitudes [9319] = 8'd119;
   assign soundFileAmplitudes [9320] = 8'd117;
   assign soundFileAmplitudes [9321] = 8'd117;
   assign soundFileAmplitudes [9322] = 8'd126;
   assign soundFileAmplitudes [9323] = 8'd136;
   assign soundFileAmplitudes [9324] = 8'd131;
   assign soundFileAmplitudes [9325] = 8'd127;
   assign soundFileAmplitudes [9326] = 8'd127;
   assign soundFileAmplitudes [9327] = 8'd129;
   assign soundFileAmplitudes [9328] = 8'd129;
   assign soundFileAmplitudes [9329] = 8'd126;
   assign soundFileAmplitudes [9330] = 8'd130;
   assign soundFileAmplitudes [9331] = 8'd142;
   assign soundFileAmplitudes [9332] = 8'd150;
   assign soundFileAmplitudes [9333] = 8'd153;
   assign soundFileAmplitudes [9334] = 8'd150;
   assign soundFileAmplitudes [9335] = 8'd152;
   assign soundFileAmplitudes [9336] = 8'd140;
   assign soundFileAmplitudes [9337] = 8'd129;
   assign soundFileAmplitudes [9338] = 8'd132;
   assign soundFileAmplitudes [9339] = 8'd135;
   assign soundFileAmplitudes [9340] = 8'd120;
   assign soundFileAmplitudes [9341] = 8'd101;
   assign soundFileAmplitudes [9342] = 8'd109;
   assign soundFileAmplitudes [9343] = 8'd114;
   assign soundFileAmplitudes [9344] = 8'd106;
   assign soundFileAmplitudes [9345] = 8'd107;
   assign soundFileAmplitudes [9346] = 8'd109;
   assign soundFileAmplitudes [9347] = 8'd112;
   assign soundFileAmplitudes [9348] = 8'd125;
   assign soundFileAmplitudes [9349] = 8'd137;
   assign soundFileAmplitudes [9350] = 8'd134;
   assign soundFileAmplitudes [9351] = 8'd118;
   assign soundFileAmplitudes [9352] = 8'd122;
   assign soundFileAmplitudes [9353] = 8'd126;
   assign soundFileAmplitudes [9354] = 8'd123;
   assign soundFileAmplitudes [9355] = 8'd124;
   assign soundFileAmplitudes [9356] = 8'd123;
   assign soundFileAmplitudes [9357] = 8'd121;
   assign soundFileAmplitudes [9358] = 8'd103;
   assign soundFileAmplitudes [9359] = 8'd97;
   assign soundFileAmplitudes [9360] = 8'd114;
   assign soundFileAmplitudes [9361] = 8'd132;
   assign soundFileAmplitudes [9362] = 8'd141;
   assign soundFileAmplitudes [9363] = 8'd142;
   assign soundFileAmplitudes [9364] = 8'd141;
   assign soundFileAmplitudes [9365] = 8'd156;
   assign soundFileAmplitudes [9366] = 8'd167;
   assign soundFileAmplitudes [9367] = 8'd158;
   assign soundFileAmplitudes [9368] = 8'd157;
   assign soundFileAmplitudes [9369] = 8'd157;
   assign soundFileAmplitudes [9370] = 8'd156;
   assign soundFileAmplitudes [9371] = 8'd128;
   assign soundFileAmplitudes [9372] = 8'd98;
   assign soundFileAmplitudes [9373] = 8'd105;
   assign soundFileAmplitudes [9374] = 8'd117;
   assign soundFileAmplitudes [9375] = 8'd111;
   assign soundFileAmplitudes [9376] = 8'd102;
   assign soundFileAmplitudes [9377] = 8'd102;
   assign soundFileAmplitudes [9378] = 8'd109;
   assign soundFileAmplitudes [9379] = 8'd120;
   assign soundFileAmplitudes [9380] = 8'd129;
   assign soundFileAmplitudes [9381] = 8'd139;
   assign soundFileAmplitudes [9382] = 8'd139;
   assign soundFileAmplitudes [9383] = 8'd136;
   assign soundFileAmplitudes [9384] = 8'd133;
   assign soundFileAmplitudes [9385] = 8'd136;
   assign soundFileAmplitudes [9386] = 8'd128;
   assign soundFileAmplitudes [9387] = 8'd113;
   assign soundFileAmplitudes [9388] = 8'd114;
   assign soundFileAmplitudes [9389] = 8'd105;
   assign soundFileAmplitudes [9390] = 8'd112;
   assign soundFileAmplitudes [9391] = 8'd126;
   assign soundFileAmplitudes [9392] = 8'd116;
   assign soundFileAmplitudes [9393] = 8'd110;
   assign soundFileAmplitudes [9394] = 8'd111;
   assign soundFileAmplitudes [9395] = 8'd121;
   assign soundFileAmplitudes [9396] = 8'd141;
   assign soundFileAmplitudes [9397] = 8'd151;
   assign soundFileAmplitudes [9398] = 8'd152;
   assign soundFileAmplitudes [9399] = 8'd150;
   assign soundFileAmplitudes [9400] = 8'd150;
   assign soundFileAmplitudes [9401] = 8'd156;
   assign soundFileAmplitudes [9402] = 8'd138;
   assign soundFileAmplitudes [9403] = 8'd123;
   assign soundFileAmplitudes [9404] = 8'd139;
   assign soundFileAmplitudes [9405] = 8'd146;
   assign soundFileAmplitudes [9406] = 8'd132;
   assign soundFileAmplitudes [9407] = 8'd110;
   assign soundFileAmplitudes [9408] = 8'd106;
   assign soundFileAmplitudes [9409] = 8'd116;
   assign soundFileAmplitudes [9410] = 8'd124;
   assign soundFileAmplitudes [9411] = 8'd127;
   assign soundFileAmplitudes [9412] = 8'd122;
   assign soundFileAmplitudes [9413] = 8'd116;
   assign soundFileAmplitudes [9414] = 8'd114;
   assign soundFileAmplitudes [9415] = 8'd112;
   assign soundFileAmplitudes [9416] = 8'd119;
   assign soundFileAmplitudes [9417] = 8'd118;
   assign soundFileAmplitudes [9418] = 8'd120;
   assign soundFileAmplitudes [9419] = 8'd111;
   assign soundFileAmplitudes [9420] = 8'd104;
   assign soundFileAmplitudes [9421] = 8'd107;
   assign soundFileAmplitudes [9422] = 8'd118;
   assign soundFileAmplitudes [9423] = 8'd134;
   assign soundFileAmplitudes [9424] = 8'd118;
   assign soundFileAmplitudes [9425] = 8'd118;
   assign soundFileAmplitudes [9426] = 8'd125;
   assign soundFileAmplitudes [9427] = 8'd133;
   assign soundFileAmplitudes [9428] = 8'd143;
   assign soundFileAmplitudes [9429] = 8'd120;
   assign soundFileAmplitudes [9430] = 8'd117;
   assign soundFileAmplitudes [9431] = 8'd143;
   assign soundFileAmplitudes [9432] = 8'd149;
   assign soundFileAmplitudes [9433] = 8'd140;
   assign soundFileAmplitudes [9434] = 8'd112;
   assign soundFileAmplitudes [9435] = 8'd113;
   assign soundFileAmplitudes [9436] = 8'd137;
   assign soundFileAmplitudes [9437] = 8'd138;
   assign soundFileAmplitudes [9438] = 8'd138;
   assign soundFileAmplitudes [9439] = 8'd140;
   assign soundFileAmplitudes [9440] = 8'd145;
   assign soundFileAmplitudes [9441] = 8'd140;
   assign soundFileAmplitudes [9442] = 8'd123;
   assign soundFileAmplitudes [9443] = 8'd117;
   assign soundFileAmplitudes [9444] = 8'd126;
   assign soundFileAmplitudes [9445] = 8'd137;
   assign soundFileAmplitudes [9446] = 8'd139;
   assign soundFileAmplitudes [9447] = 8'd125;
   assign soundFileAmplitudes [9448] = 8'd116;
   assign soundFileAmplitudes [9449] = 8'd113;
   assign soundFileAmplitudes [9450] = 8'd105;
   assign soundFileAmplitudes [9451] = 8'd118;
   assign soundFileAmplitudes [9452] = 8'd124;
   assign soundFileAmplitudes [9453] = 8'd132;
   assign soundFileAmplitudes [9454] = 8'd135;
   assign soundFileAmplitudes [9455] = 8'd126;
   assign soundFileAmplitudes [9456] = 8'd109;
   assign soundFileAmplitudes [9457] = 8'd101;
   assign soundFileAmplitudes [9458] = 8'd115;
   assign soundFileAmplitudes [9459] = 8'd118;
   assign soundFileAmplitudes [9460] = 8'd116;
   assign soundFileAmplitudes [9461] = 8'd102;
   assign soundFileAmplitudes [9462] = 8'd120;
   assign soundFileAmplitudes [9463] = 8'd137;
   assign soundFileAmplitudes [9464] = 8'd132;
   assign soundFileAmplitudes [9465] = 8'd105;
   assign soundFileAmplitudes [9466] = 8'd104;
   assign soundFileAmplitudes [9467] = 8'd136;
   assign soundFileAmplitudes [9468] = 8'd142;
   assign soundFileAmplitudes [9469] = 8'd139;
   assign soundFileAmplitudes [9470] = 8'd142;
   assign soundFileAmplitudes [9471] = 8'd158;
   assign soundFileAmplitudes [9472] = 8'd159;
   assign soundFileAmplitudes [9473] = 8'd155;
   assign soundFileAmplitudes [9474] = 8'd145;
   assign soundFileAmplitudes [9475] = 8'd138;
   assign soundFileAmplitudes [9476] = 8'd120;
   assign soundFileAmplitudes [9477] = 8'd108;
   assign soundFileAmplitudes [9478] = 8'd112;
   assign soundFileAmplitudes [9479] = 8'd115;
   assign soundFileAmplitudes [9480] = 8'd107;
   assign soundFileAmplitudes [9481] = 8'd106;
   assign soundFileAmplitudes [9482] = 8'd125;
   assign soundFileAmplitudes [9483] = 8'd133;
   assign soundFileAmplitudes [9484] = 8'd136;
   assign soundFileAmplitudes [9485] = 8'd136;
   assign soundFileAmplitudes [9486] = 8'd137;
   assign soundFileAmplitudes [9487] = 8'd134;
   assign soundFileAmplitudes [9488] = 8'd133;
   assign soundFileAmplitudes [9489] = 8'd130;
   assign soundFileAmplitudes [9490] = 8'd135;
   assign soundFileAmplitudes [9491] = 8'd110;
   assign soundFileAmplitudes [9492] = 8'd93;
   assign soundFileAmplitudes [9493] = 8'd99;
   assign soundFileAmplitudes [9494] = 8'd101;
   assign soundFileAmplitudes [9495] = 8'd100;
   assign soundFileAmplitudes [9496] = 8'd85;
   assign soundFileAmplitudes [9497] = 8'd106;
   assign soundFileAmplitudes [9498] = 8'd129;
   assign soundFileAmplitudes [9499] = 8'd134;
   assign soundFileAmplitudes [9500] = 8'd131;
   assign soundFileAmplitudes [9501] = 8'd138;
   assign soundFileAmplitudes [9502] = 8'd160;
   assign soundFileAmplitudes [9503] = 8'd168;
   assign soundFileAmplitudes [9504] = 8'd166;
   assign soundFileAmplitudes [9505] = 8'd170;
   assign soundFileAmplitudes [9506] = 8'd159;
   assign soundFileAmplitudes [9507] = 8'd145;
   assign soundFileAmplitudes [9508] = 8'd133;
   assign soundFileAmplitudes [9509] = 8'd120;
   assign soundFileAmplitudes [9510] = 8'd113;
   assign soundFileAmplitudes [9511] = 8'd95;
   assign soundFileAmplitudes [9512] = 8'd100;
   assign soundFileAmplitudes [9513] = 8'd116;
   assign soundFileAmplitudes [9514] = 8'd124;
   assign soundFileAmplitudes [9515] = 8'd131;
   assign soundFileAmplitudes [9516] = 8'd129;
   assign soundFileAmplitudes [9517] = 8'd131;
   assign soundFileAmplitudes [9518] = 8'd136;
   assign soundFileAmplitudes [9519] = 8'd135;
   assign soundFileAmplitudes [9520] = 8'd143;
   assign soundFileAmplitudes [9521] = 8'd141;
   assign soundFileAmplitudes [9522] = 8'd122;
   assign soundFileAmplitudes [9523] = 8'd125;
   assign soundFileAmplitudes [9524] = 8'd131;
   assign soundFileAmplitudes [9525] = 8'd128;
   assign soundFileAmplitudes [9526] = 8'd93;
   assign soundFileAmplitudes [9527] = 8'd65;
   assign soundFileAmplitudes [9528] = 8'd79;
   assign soundFileAmplitudes [9529] = 8'd89;
   assign soundFileAmplitudes [9530] = 8'd103;
   assign soundFileAmplitudes [9531] = 8'd121;
   assign soundFileAmplitudes [9532] = 8'd131;
   assign soundFileAmplitudes [9533] = 8'd136;
   assign soundFileAmplitudes [9534] = 8'd145;
   assign soundFileAmplitudes [9535] = 8'd149;
   assign soundFileAmplitudes [9536] = 8'd160;
   assign soundFileAmplitudes [9537] = 8'd164;
   assign soundFileAmplitudes [9538] = 8'd153;
   assign soundFileAmplitudes [9539] = 8'd141;
   assign soundFileAmplitudes [9540] = 8'd142;
   assign soundFileAmplitudes [9541] = 8'd134;
   assign soundFileAmplitudes [9542] = 8'd124;
   assign soundFileAmplitudes [9543] = 8'd135;
   assign soundFileAmplitudes [9544] = 8'd129;
   assign soundFileAmplitudes [9545] = 8'd123;
   assign soundFileAmplitudes [9546] = 8'd118;
   assign soundFileAmplitudes [9547] = 8'd116;
   assign soundFileAmplitudes [9548] = 8'd119;
   assign soundFileAmplitudes [9549] = 8'd123;
   assign soundFileAmplitudes [9550] = 8'd131;
   assign soundFileAmplitudes [9551] = 8'd126;
   assign soundFileAmplitudes [9552] = 8'd113;
   assign soundFileAmplitudes [9553] = 8'd108;
   assign soundFileAmplitudes [9554] = 8'd115;
   assign soundFileAmplitudes [9555] = 8'd130;
   assign soundFileAmplitudes [9556] = 8'd121;
   assign soundFileAmplitudes [9557] = 8'd98;
   assign soundFileAmplitudes [9558] = 8'd108;
   assign soundFileAmplitudes [9559] = 8'd124;
   assign soundFileAmplitudes [9560] = 8'd121;
   assign soundFileAmplitudes [9561] = 8'd109;
   assign soundFileAmplitudes [9562] = 8'd118;
   assign soundFileAmplitudes [9563] = 8'd130;
   assign soundFileAmplitudes [9564] = 8'd132;
   assign soundFileAmplitudes [9565] = 8'd134;
   assign soundFileAmplitudes [9566] = 8'd131;
   assign soundFileAmplitudes [9567] = 8'd137;
   assign soundFileAmplitudes [9568] = 8'd140;
   assign soundFileAmplitudes [9569] = 8'd137;
   assign soundFileAmplitudes [9570] = 8'd140;
   assign soundFileAmplitudes [9571] = 8'd138;
   assign soundFileAmplitudes [9572] = 8'd137;
   assign soundFileAmplitudes [9573] = 8'd143;
   assign soundFileAmplitudes [9574] = 8'd142;
   assign soundFileAmplitudes [9575] = 8'd139;
   assign soundFileAmplitudes [9576] = 8'd127;
   assign soundFileAmplitudes [9577] = 8'd125;
   assign soundFileAmplitudes [9578] = 8'd132;
   assign soundFileAmplitudes [9579] = 8'd128;
   assign soundFileAmplitudes [9580] = 8'd121;
   assign soundFileAmplitudes [9581] = 8'd118;
   assign soundFileAmplitudes [9582] = 8'd109;
   assign soundFileAmplitudes [9583] = 8'd105;
   assign soundFileAmplitudes [9584] = 8'd99;
   assign soundFileAmplitudes [9585] = 8'd103;
   assign soundFileAmplitudes [9586] = 8'd123;
   assign soundFileAmplitudes [9587] = 8'd113;
   assign soundFileAmplitudes [9588] = 8'd97;
   assign soundFileAmplitudes [9589] = 8'd92;
   assign soundFileAmplitudes [9590] = 8'd113;
   assign soundFileAmplitudes [9591] = 8'd124;
   assign soundFileAmplitudes [9592] = 8'd122;
   assign soundFileAmplitudes [9593] = 8'd122;
   assign soundFileAmplitudes [9594] = 8'd128;
   assign soundFileAmplitudes [9595] = 8'd148;
   assign soundFileAmplitudes [9596] = 8'd151;
   assign soundFileAmplitudes [9597] = 8'd139;
   assign soundFileAmplitudes [9598] = 8'd131;
   assign soundFileAmplitudes [9599] = 8'd138;
   assign soundFileAmplitudes [9600] = 8'd143;
   assign soundFileAmplitudes [9601] = 8'd139;
   assign soundFileAmplitudes [9602] = 8'd126;
   assign soundFileAmplitudes [9603] = 8'd112;
   assign soundFileAmplitudes [9604] = 8'd117;
   assign soundFileAmplitudes [9605] = 8'd137;
   assign soundFileAmplitudes [9606] = 8'd150;
   assign soundFileAmplitudes [9607] = 8'd155;
   assign soundFileAmplitudes [9608] = 8'd149;
   assign soundFileAmplitudes [9609] = 8'd138;
   assign soundFileAmplitudes [9610] = 8'd134;
   assign soundFileAmplitudes [9611] = 8'd126;
   assign soundFileAmplitudes [9612] = 8'd133;
   assign soundFileAmplitudes [9613] = 8'd140;
   assign soundFileAmplitudes [9614] = 8'd129;
   assign soundFileAmplitudes [9615] = 8'd108;
   assign soundFileAmplitudes [9616] = 8'd99;
   assign soundFileAmplitudes [9617] = 8'd106;
   assign soundFileAmplitudes [9618] = 8'd103;
   assign soundFileAmplitudes [9619] = 8'd97;
   assign soundFileAmplitudes [9620] = 8'd99;
   assign soundFileAmplitudes [9621] = 8'd113;
   assign soundFileAmplitudes [9622] = 8'd118;
   assign soundFileAmplitudes [9623] = 8'd125;
   assign soundFileAmplitudes [9624] = 8'd140;
   assign soundFileAmplitudes [9625] = 8'd145;
   assign soundFileAmplitudes [9626] = 8'd146;
   assign soundFileAmplitudes [9627] = 8'd140;
   assign soundFileAmplitudes [9628] = 8'd142;
   assign soundFileAmplitudes [9629] = 8'd143;
   assign soundFileAmplitudes [9630] = 8'd137;
   assign soundFileAmplitudes [9631] = 8'd123;
   assign soundFileAmplitudes [9632] = 8'd113;
   assign soundFileAmplitudes [9633] = 8'd104;
   assign soundFileAmplitudes [9634] = 8'd99;
   assign soundFileAmplitudes [9635] = 8'd109;
   assign soundFileAmplitudes [9636] = 8'd119;
   assign soundFileAmplitudes [9637] = 8'd127;
   assign soundFileAmplitudes [9638] = 8'd128;
   assign soundFileAmplitudes [9639] = 8'd129;
   assign soundFileAmplitudes [9640] = 8'd133;
   assign soundFileAmplitudes [9641] = 8'd148;
   assign soundFileAmplitudes [9642] = 8'd164;
   assign soundFileAmplitudes [9643] = 8'd168;
   assign soundFileAmplitudes [9644] = 8'd146;
   assign soundFileAmplitudes [9645] = 8'd138;
   assign soundFileAmplitudes [9646] = 8'd145;
   assign soundFileAmplitudes [9647] = 8'd141;
   assign soundFileAmplitudes [9648] = 8'd126;
   assign soundFileAmplitudes [9649] = 8'd93;
   assign soundFileAmplitudes [9650] = 8'd80;
   assign soundFileAmplitudes [9651] = 8'd91;
   assign soundFileAmplitudes [9652] = 8'd95;
   assign soundFileAmplitudes [9653] = 8'd99;
   assign soundFileAmplitudes [9654] = 8'd114;
   assign soundFileAmplitudes [9655] = 8'd132;
   assign soundFileAmplitudes [9656] = 8'd138;
   assign soundFileAmplitudes [9657] = 8'd137;
   assign soundFileAmplitudes [9658] = 8'd139;
   assign soundFileAmplitudes [9659] = 8'd135;
   assign soundFileAmplitudes [9660] = 8'd146;
   assign soundFileAmplitudes [9661] = 8'd141;
   assign soundFileAmplitudes [9662] = 8'd134;
   assign soundFileAmplitudes [9663] = 8'd125;
   assign soundFileAmplitudes [9664] = 8'd120;
   assign soundFileAmplitudes [9665] = 8'd120;
   assign soundFileAmplitudes [9666] = 8'd108;
   assign soundFileAmplitudes [9667] = 8'd110;
   assign soundFileAmplitudes [9668] = 8'd103;
   assign soundFileAmplitudes [9669] = 8'd108;
   assign soundFileAmplitudes [9670] = 8'd124;
   assign soundFileAmplitudes [9671] = 8'd133;
   assign soundFileAmplitudes [9672] = 8'd141;
   assign soundFileAmplitudes [9673] = 8'd134;
   assign soundFileAmplitudes [9674] = 8'd128;
   assign soundFileAmplitudes [9675] = 8'd143;
   assign soundFileAmplitudes [9676] = 8'd146;
   assign soundFileAmplitudes [9677] = 8'd151;
   assign soundFileAmplitudes [9678] = 8'd138;
   assign soundFileAmplitudes [9679] = 8'd122;
   assign soundFileAmplitudes [9680] = 8'd136;
   assign soundFileAmplitudes [9681] = 8'd138;
   assign soundFileAmplitudes [9682] = 8'd132;
   assign soundFileAmplitudes [9683] = 8'd123;
   assign soundFileAmplitudes [9684] = 8'd113;
   assign soundFileAmplitudes [9685] = 8'd108;
   assign soundFileAmplitudes [9686] = 8'd111;
   assign soundFileAmplitudes [9687] = 8'd114;
   assign soundFileAmplitudes [9688] = 8'd119;
   assign soundFileAmplitudes [9689] = 8'd128;
   assign soundFileAmplitudes [9690] = 8'd130;
   assign soundFileAmplitudes [9691] = 8'd124;
   assign soundFileAmplitudes [9692] = 8'd111;
   assign soundFileAmplitudes [9693] = 8'd107;
   assign soundFileAmplitudes [9694] = 8'd116;
   assign soundFileAmplitudes [9695] = 8'd121;
   assign soundFileAmplitudes [9696] = 8'd135;
   assign soundFileAmplitudes [9697] = 8'd143;
   assign soundFileAmplitudes [9698] = 8'd143;
   assign soundFileAmplitudes [9699] = 8'd134;
   assign soundFileAmplitudes [9700] = 8'd108;
   assign soundFileAmplitudes [9701] = 8'd112;
   assign soundFileAmplitudes [9702] = 8'd115;
   assign soundFileAmplitudes [9703] = 8'd124;
   assign soundFileAmplitudes [9704] = 8'd131;
   assign soundFileAmplitudes [9705] = 8'd116;
   assign soundFileAmplitudes [9706] = 8'd116;
   assign soundFileAmplitudes [9707] = 8'd113;
   assign soundFileAmplitudes [9708] = 8'd119;
   assign soundFileAmplitudes [9709] = 8'd124;
   assign soundFileAmplitudes [9710] = 8'd125;
   assign soundFileAmplitudes [9711] = 8'd149;
   assign soundFileAmplitudes [9712] = 8'd156;
   assign soundFileAmplitudes [9713] = 8'd146;
   assign soundFileAmplitudes [9714] = 8'd139;
   assign soundFileAmplitudes [9715] = 8'd144;
   assign soundFileAmplitudes [9716] = 8'd151;
   assign soundFileAmplitudes [9717] = 8'd149;
   assign soundFileAmplitudes [9718] = 8'd138;
   assign soundFileAmplitudes [9719] = 8'd121;
   assign soundFileAmplitudes [9720] = 8'd108;
   assign soundFileAmplitudes [9721] = 8'd100;
   assign soundFileAmplitudes [9722] = 8'd101;
   assign soundFileAmplitudes [9723] = 8'd106;
   assign soundFileAmplitudes [9724] = 8'd118;
   assign soundFileAmplitudes [9725] = 8'd105;
   assign soundFileAmplitudes [9726] = 8'd97;
   assign soundFileAmplitudes [9727] = 8'd107;
   assign soundFileAmplitudes [9728] = 8'd122;
   assign soundFileAmplitudes [9729] = 8'd142;
   assign soundFileAmplitudes [9730] = 8'd143;
   assign soundFileAmplitudes [9731] = 8'd146;
   assign soundFileAmplitudes [9732] = 8'd145;
   assign soundFileAmplitudes [9733] = 8'd144;
   assign soundFileAmplitudes [9734] = 8'd137;
   assign soundFileAmplitudes [9735] = 8'd128;
   assign soundFileAmplitudes [9736] = 8'd125;
   assign soundFileAmplitudes [9737] = 8'd120;
   assign soundFileAmplitudes [9738] = 8'd110;
   assign soundFileAmplitudes [9739] = 8'd112;
   assign soundFileAmplitudes [9740] = 8'd114;
   assign soundFileAmplitudes [9741] = 8'd102;
   assign soundFileAmplitudes [9742] = 8'd107;
   assign soundFileAmplitudes [9743] = 8'd121;
   assign soundFileAmplitudes [9744] = 8'd130;
   assign soundFileAmplitudes [9745] = 8'd142;
   assign soundFileAmplitudes [9746] = 8'd154;
   assign soundFileAmplitudes [9747] = 8'd156;
   assign soundFileAmplitudes [9748] = 8'd153;
   assign soundFileAmplitudes [9749] = 8'd141;
   assign soundFileAmplitudes [9750] = 8'd135;
   assign soundFileAmplitudes [9751] = 8'd138;
   assign soundFileAmplitudes [9752] = 8'd136;
   assign soundFileAmplitudes [9753] = 8'd126;
   assign soundFileAmplitudes [9754] = 8'd116;
   assign soundFileAmplitudes [9755] = 8'd105;
   assign soundFileAmplitudes [9756] = 8'd101;
   assign soundFileAmplitudes [9757] = 8'd101;
   assign soundFileAmplitudes [9758] = 8'd109;
   assign soundFileAmplitudes [9759] = 8'd113;
   assign soundFileAmplitudes [9760] = 8'd116;
   assign soundFileAmplitudes [9761] = 8'd118;
   assign soundFileAmplitudes [9762] = 8'd115;
   assign soundFileAmplitudes [9763] = 8'd126;
   assign soundFileAmplitudes [9764] = 8'd132;
   assign soundFileAmplitudes [9765] = 8'd144;
   assign soundFileAmplitudes [9766] = 8'd145;
   assign soundFileAmplitudes [9767] = 8'd137;
   assign soundFileAmplitudes [9768] = 8'd122;
   assign soundFileAmplitudes [9769] = 8'd120;
   assign soundFileAmplitudes [9770] = 8'd136;
   assign soundFileAmplitudes [9771] = 8'd138;
   assign soundFileAmplitudes [9772] = 8'd115;
   assign soundFileAmplitudes [9773] = 8'd101;
   assign soundFileAmplitudes [9774] = 8'd116;
   assign soundFileAmplitudes [9775] = 8'd136;
   assign soundFileAmplitudes [9776] = 8'd145;
   assign soundFileAmplitudes [9777] = 8'd132;
   assign soundFileAmplitudes [9778] = 8'd129;
   assign soundFileAmplitudes [9779] = 8'd133;
   assign soundFileAmplitudes [9780] = 8'd145;
   assign soundFileAmplitudes [9781] = 8'd148;
   assign soundFileAmplitudes [9782] = 8'd139;
   assign soundFileAmplitudes [9783] = 8'd136;
   assign soundFileAmplitudes [9784] = 8'd128;
   assign soundFileAmplitudes [9785] = 8'd124;
   assign soundFileAmplitudes [9786] = 8'd129;
   assign soundFileAmplitudes [9787] = 8'd119;
   assign soundFileAmplitudes [9788] = 8'd108;
   assign soundFileAmplitudes [9789] = 8'd113;
   assign soundFileAmplitudes [9790] = 8'd125;
   assign soundFileAmplitudes [9791] = 8'd136;
   assign soundFileAmplitudes [9792] = 8'd138;
   assign soundFileAmplitudes [9793] = 8'd135;
   assign soundFileAmplitudes [9794] = 8'd122;
   assign soundFileAmplitudes [9795] = 8'd116;
   assign soundFileAmplitudes [9796] = 8'd117;
   assign soundFileAmplitudes [9797] = 8'd136;
   assign soundFileAmplitudes [9798] = 8'd135;
   assign soundFileAmplitudes [9799] = 8'd129;
   assign soundFileAmplitudes [9800] = 8'd124;
   assign soundFileAmplitudes [9801] = 8'd117;
   assign soundFileAmplitudes [9802] = 8'd100;
   assign soundFileAmplitudes [9803] = 8'd73;
   assign soundFileAmplitudes [9804] = 8'd91;
   assign soundFileAmplitudes [9805] = 8'd104;
   assign soundFileAmplitudes [9806] = 8'd123;
   assign soundFileAmplitudes [9807] = 8'd134;
   assign soundFileAmplitudes [9808] = 8'd137;
   assign soundFileAmplitudes [9809] = 8'd143;
   assign soundFileAmplitudes [9810] = 8'd144;
   assign soundFileAmplitudes [9811] = 8'd152;
   assign soundFileAmplitudes [9812] = 8'd148;
   assign soundFileAmplitudes [9813] = 8'd149;
   assign soundFileAmplitudes [9814] = 8'd155;
   assign soundFileAmplitudes [9815] = 8'd144;
   assign soundFileAmplitudes [9816] = 8'd127;
   assign soundFileAmplitudes [9817] = 8'd127;
   assign soundFileAmplitudes [9818] = 8'd134;
   assign soundFileAmplitudes [9819] = 8'd126;
   assign soundFileAmplitudes [9820] = 8'd120;
   assign soundFileAmplitudes [9821] = 8'd121;
   assign soundFileAmplitudes [9822] = 8'd117;
   assign soundFileAmplitudes [9823] = 8'd115;
   assign soundFileAmplitudes [9824] = 8'd116;
   assign soundFileAmplitudes [9825] = 8'd129;
   assign soundFileAmplitudes [9826] = 8'd133;
   assign soundFileAmplitudes [9827] = 8'd131;
   assign soundFileAmplitudes [9828] = 8'd126;
   assign soundFileAmplitudes [9829] = 8'd121;
   assign soundFileAmplitudes [9830] = 8'd116;
   assign soundFileAmplitudes [9831] = 8'd105;
   assign soundFileAmplitudes [9832] = 8'd104;
   assign soundFileAmplitudes [9833] = 8'd101;
   assign soundFileAmplitudes [9834] = 8'd109;
   assign soundFileAmplitudes [9835] = 8'd117;
   assign soundFileAmplitudes [9836] = 8'd120;
   assign soundFileAmplitudes [9837] = 8'd108;
   assign soundFileAmplitudes [9838] = 8'd97;
   assign soundFileAmplitudes [9839] = 8'd117;
   assign soundFileAmplitudes [9840] = 8'd134;
   assign soundFileAmplitudes [9841] = 8'd144;
   assign soundFileAmplitudes [9842] = 8'd153;
   assign soundFileAmplitudes [9843] = 8'd151;
   assign soundFileAmplitudes [9844] = 8'd144;
   assign soundFileAmplitudes [9845] = 8'd147;
   assign soundFileAmplitudes [9846] = 8'd147;
   assign soundFileAmplitudes [9847] = 8'd144;
   assign soundFileAmplitudes [9848] = 8'd140;
   assign soundFileAmplitudes [9849] = 8'd131;
   assign soundFileAmplitudes [9850] = 8'd117;
   assign soundFileAmplitudes [9851] = 8'd118;
   assign soundFileAmplitudes [9852] = 8'd122;
   assign soundFileAmplitudes [9853] = 8'd117;
   assign soundFileAmplitudes [9854] = 8'd121;
   assign soundFileAmplitudes [9855] = 8'd118;
   assign soundFileAmplitudes [9856] = 8'd121;
   assign soundFileAmplitudes [9857] = 8'd124;
   assign soundFileAmplitudes [9858] = 8'd114;
   assign soundFileAmplitudes [9859] = 8'd119;
   assign soundFileAmplitudes [9860] = 8'd130;
   assign soundFileAmplitudes [9861] = 8'd128;
   assign soundFileAmplitudes [9862] = 8'd119;
   assign soundFileAmplitudes [9863] = 8'd115;
   assign soundFileAmplitudes [9864] = 8'd121;
   assign soundFileAmplitudes [9865] = 8'd129;
   assign soundFileAmplitudes [9866] = 8'd123;
   assign soundFileAmplitudes [9867] = 8'd118;
   assign soundFileAmplitudes [9868] = 8'd114;
   assign soundFileAmplitudes [9869] = 8'd111;
   assign soundFileAmplitudes [9870] = 8'd133;
   assign soundFileAmplitudes [9871] = 8'd148;
   assign soundFileAmplitudes [9872] = 8'd144;
   assign soundFileAmplitudes [9873] = 8'd123;
   assign soundFileAmplitudes [9874] = 8'd113;
   assign soundFileAmplitudes [9875] = 8'd105;
   assign soundFileAmplitudes [9876] = 8'd121;
   assign soundFileAmplitudes [9877] = 8'd135;
   assign soundFileAmplitudes [9878] = 8'd136;
   assign soundFileAmplitudes [9879] = 8'd138;
   assign soundFileAmplitudes [9880] = 8'd111;
   assign soundFileAmplitudes [9881] = 8'd101;
   assign soundFileAmplitudes [9882] = 8'd116;
   assign soundFileAmplitudes [9883] = 8'd137;
   assign soundFileAmplitudes [9884] = 8'd147;
   assign soundFileAmplitudes [9885] = 8'd143;
   assign soundFileAmplitudes [9886] = 8'd134;
   assign soundFileAmplitudes [9887] = 8'd142;
   assign soundFileAmplitudes [9888] = 8'd136;
   assign soundFileAmplitudes [9889] = 8'd129;
   assign soundFileAmplitudes [9890] = 8'd136;
   assign soundFileAmplitudes [9891] = 8'd128;
   assign soundFileAmplitudes [9892] = 8'd120;
   assign soundFileAmplitudes [9893] = 8'd103;
   assign soundFileAmplitudes [9894] = 8'd105;
   assign soundFileAmplitudes [9895] = 8'd125;
   assign soundFileAmplitudes [9896] = 8'd137;
   assign soundFileAmplitudes [9897] = 8'd134;
   assign soundFileAmplitudes [9898] = 8'd121;
   assign soundFileAmplitudes [9899] = 8'd113;
   assign soundFileAmplitudes [9900] = 8'd117;
   assign soundFileAmplitudes [9901] = 8'd116;
   assign soundFileAmplitudes [9902] = 8'd131;
   assign soundFileAmplitudes [9903] = 8'd144;
   assign soundFileAmplitudes [9904] = 8'd142;
   assign soundFileAmplitudes [9905] = 8'd137;
   assign soundFileAmplitudes [9906] = 8'd144;
   assign soundFileAmplitudes [9907] = 8'd142;
   assign soundFileAmplitudes [9908] = 8'd126;
   assign soundFileAmplitudes [9909] = 8'd113;
   assign soundFileAmplitudes [9910] = 8'd101;
   assign soundFileAmplitudes [9911] = 8'd98;
   assign soundFileAmplitudes [9912] = 8'd101;
   assign soundFileAmplitudes [9913] = 8'd117;
   assign soundFileAmplitudes [9914] = 8'd122;
   assign soundFileAmplitudes [9915] = 8'd120;
   assign soundFileAmplitudes [9916] = 8'd120;
   assign soundFileAmplitudes [9917] = 8'd127;
   assign soundFileAmplitudes [9918] = 8'd147;
   assign soundFileAmplitudes [9919] = 8'd163;
   assign soundFileAmplitudes [9920] = 8'd152;
   assign soundFileAmplitudes [9921] = 8'd137;
   assign soundFileAmplitudes [9922] = 8'd141;
   assign soundFileAmplitudes [9923] = 8'd147;
   assign soundFileAmplitudes [9924] = 8'd146;
   assign soundFileAmplitudes [9925] = 8'd130;
   assign soundFileAmplitudes [9926] = 8'd129;
   assign soundFileAmplitudes [9927] = 8'd128;
   assign soundFileAmplitudes [9928] = 8'd126;
   assign soundFileAmplitudes [9929] = 8'd118;
   assign soundFileAmplitudes [9930] = 8'd106;
   assign soundFileAmplitudes [9931] = 8'd116;
   assign soundFileAmplitudes [9932] = 8'd121;
   assign soundFileAmplitudes [9933] = 8'd134;
   assign soundFileAmplitudes [9934] = 8'd139;
   assign soundFileAmplitudes [9935] = 8'd131;
   assign soundFileAmplitudes [9936] = 8'd131;
   assign soundFileAmplitudes [9937] = 8'd132;
   assign soundFileAmplitudes [9938] = 8'd129;
   assign soundFileAmplitudes [9939] = 8'd121;
   assign soundFileAmplitudes [9940] = 8'd127;
   assign soundFileAmplitudes [9941] = 8'd123;
   assign soundFileAmplitudes [9942] = 8'd107;
   assign soundFileAmplitudes [9943] = 8'd92;
   assign soundFileAmplitudes [9944] = 8'd91;
   assign soundFileAmplitudes [9945] = 8'd105;
   assign soundFileAmplitudes [9946] = 8'd116;
   assign soundFileAmplitudes [9947] = 8'd123;
   assign soundFileAmplitudes [9948] = 8'd126;
   assign soundFileAmplitudes [9949] = 8'd127;
   assign soundFileAmplitudes [9950] = 8'd114;
   assign soundFileAmplitudes [9951] = 8'd116;
   assign soundFileAmplitudes [9952] = 8'd123;
   assign soundFileAmplitudes [9953] = 8'd141;
   assign soundFileAmplitudes [9954] = 8'd158;
   assign soundFileAmplitudes [9955] = 8'd142;
   assign soundFileAmplitudes [9956] = 8'd118;
   assign soundFileAmplitudes [9957] = 8'd116;
   assign soundFileAmplitudes [9958] = 8'd122;
   assign soundFileAmplitudes [9959] = 8'd125;
   assign soundFileAmplitudes [9960] = 8'd129;
   assign soundFileAmplitudes [9961] = 8'd124;
   assign soundFileAmplitudes [9962] = 8'd122;
   assign soundFileAmplitudes [9963] = 8'd126;
   assign soundFileAmplitudes [9964] = 8'd142;
   assign soundFileAmplitudes [9965] = 8'd153;
   assign soundFileAmplitudes [9966] = 8'd160;
   assign soundFileAmplitudes [9967] = 8'd162;
   assign soundFileAmplitudes [9968] = 8'd149;
   assign soundFileAmplitudes [9969] = 8'd141;
   assign soundFileAmplitudes [9970] = 8'd130;
   assign soundFileAmplitudes [9971] = 8'd123;
   assign soundFileAmplitudes [9972] = 8'd116;
   assign soundFileAmplitudes [9973] = 8'd99;
   assign soundFileAmplitudes [9974] = 8'd92;
   assign soundFileAmplitudes [9975] = 8'd99;
   assign soundFileAmplitudes [9976] = 8'd109;
   assign soundFileAmplitudes [9977] = 8'd111;
   assign soundFileAmplitudes [9978] = 8'd95;
   assign soundFileAmplitudes [9979] = 8'd93;
   assign soundFileAmplitudes [9980] = 8'd114;
   assign soundFileAmplitudes [9981] = 8'd124;
   assign soundFileAmplitudes [9982] = 8'd125;
   assign soundFileAmplitudes [9983] = 8'd137;
   assign soundFileAmplitudes [9984] = 8'd145;
   assign soundFileAmplitudes [9985] = 8'd145;
   assign soundFileAmplitudes [9986] = 8'd137;
   assign soundFileAmplitudes [9987] = 8'd123;
   assign soundFileAmplitudes [9988] = 8'd129;
   assign soundFileAmplitudes [9989] = 8'd136;
   assign soundFileAmplitudes [9990] = 8'd128;
   assign soundFileAmplitudes [9991] = 8'd115;
   assign soundFileAmplitudes [9992] = 8'd113;
   assign soundFileAmplitudes [9993] = 8'd117;
   assign soundFileAmplitudes [9994] = 8'd124;
   assign soundFileAmplitudes [9995] = 8'd142;
   assign soundFileAmplitudes [9996] = 8'd147;
   assign soundFileAmplitudes [9997] = 8'd148;
   assign soundFileAmplitudes [9998] = 8'd158;
   assign soundFileAmplitudes [9999] = 8'd165;
   assign soundFileAmplitudes [10000] = 8'd156;
   assign soundFileAmplitudes [10001] = 8'd140;
   assign soundFileAmplitudes [10002] = 8'd144;
   assign soundFileAmplitudes [10003] = 8'd127;
   assign soundFileAmplitudes [10004] = 8'd110;
   assign soundFileAmplitudes [10005] = 8'd98;
   assign soundFileAmplitudes [10006] = 8'd92;
   assign soundFileAmplitudes [10007] = 8'd103;
   assign soundFileAmplitudes [10008] = 8'd103;
   assign soundFileAmplitudes [10009] = 8'd99;
   assign soundFileAmplitudes [10010] = 8'd101;
   assign soundFileAmplitudes [10011] = 8'd110;
   assign soundFileAmplitudes [10012] = 8'd122;
   assign soundFileAmplitudes [10013] = 8'd115;
   assign soundFileAmplitudes [10014] = 8'd100;
   assign soundFileAmplitudes [10015] = 8'd106;
   assign soundFileAmplitudes [10016] = 8'd128;
   assign soundFileAmplitudes [10017] = 8'd139;
   assign soundFileAmplitudes [10018] = 8'd123;
   assign soundFileAmplitudes [10019] = 8'd123;
   assign soundFileAmplitudes [10020] = 8'd111;
   assign soundFileAmplitudes [10021] = 8'd114;
   assign soundFileAmplitudes [10022] = 8'd122;
   assign soundFileAmplitudes [10023] = 8'd124;
   assign soundFileAmplitudes [10024] = 8'd134;
   assign soundFileAmplitudes [10025] = 8'd142;
   assign soundFileAmplitudes [10026] = 8'd139;
   assign soundFileAmplitudes [10027] = 8'd140;
   assign soundFileAmplitudes [10028] = 8'd158;
   assign soundFileAmplitudes [10029] = 8'd160;
   assign soundFileAmplitudes [10030] = 8'd166;
   assign soundFileAmplitudes [10031] = 8'd161;
   assign soundFileAmplitudes [10032] = 8'd150;
   assign soundFileAmplitudes [10033] = 8'd144;
   assign soundFileAmplitudes [10034] = 8'd136;
   assign soundFileAmplitudes [10035] = 8'd116;
   assign soundFileAmplitudes [10036] = 8'd111;
   assign soundFileAmplitudes [10037] = 8'd125;
   assign soundFileAmplitudes [10038] = 8'd127;
   assign soundFileAmplitudes [10039] = 8'd115;
   assign soundFileAmplitudes [10040] = 8'd102;
   assign soundFileAmplitudes [10041] = 8'd93;
   assign soundFileAmplitudes [10042] = 8'd101;
   assign soundFileAmplitudes [10043] = 8'd111;
   assign soundFileAmplitudes [10044] = 8'd115;
   assign soundFileAmplitudes [10045] = 8'd122;
   assign soundFileAmplitudes [10046] = 8'd137;
   assign soundFileAmplitudes [10047] = 8'd149;
   assign soundFileAmplitudes [10048] = 8'd135;
   assign soundFileAmplitudes [10049] = 8'd110;
   assign soundFileAmplitudes [10050] = 8'd109;
   assign soundFileAmplitudes [10051] = 8'd117;
   assign soundFileAmplitudes [10052] = 8'd114;
   assign soundFileAmplitudes [10053] = 8'd114;
   assign soundFileAmplitudes [10054] = 8'd111;
   assign soundFileAmplitudes [10055] = 8'd114;
   assign soundFileAmplitudes [10056] = 8'd117;
   assign soundFileAmplitudes [10057] = 8'd133;
   assign soundFileAmplitudes [10058] = 8'd142;
   assign soundFileAmplitudes [10059] = 8'd137;
   assign soundFileAmplitudes [10060] = 8'd144;
   assign soundFileAmplitudes [10061] = 8'd158;
   assign soundFileAmplitudes [10062] = 8'd165;
   assign soundFileAmplitudes [10063] = 8'd170;
   assign soundFileAmplitudes [10064] = 8'd166;
   assign soundFileAmplitudes [10065] = 8'd153;
   assign soundFileAmplitudes [10066] = 8'd129;
   assign soundFileAmplitudes [10067] = 8'd111;
   assign soundFileAmplitudes [10068] = 8'd118;
   assign soundFileAmplitudes [10069] = 8'd129;
   assign soundFileAmplitudes [10070] = 8'd128;
   assign soundFileAmplitudes [10071] = 8'd113;
   assign soundFileAmplitudes [10072] = 8'd105;
   assign soundFileAmplitudes [10073] = 8'd106;
   assign soundFileAmplitudes [10074] = 8'd104;
   assign soundFileAmplitudes [10075] = 8'd103;
   assign soundFileAmplitudes [10076] = 8'd100;
   assign soundFileAmplitudes [10077] = 8'd103;
   assign soundFileAmplitudes [10078] = 8'd123;
   assign soundFileAmplitudes [10079] = 8'd122;
   assign soundFileAmplitudes [10080] = 8'd112;
   assign soundFileAmplitudes [10081] = 8'd110;
   assign soundFileAmplitudes [10082] = 8'd120;
   assign soundFileAmplitudes [10083] = 8'd134;
   assign soundFileAmplitudes [10084] = 8'd130;
   assign soundFileAmplitudes [10085] = 8'd114;
   assign soundFileAmplitudes [10086] = 8'd109;
   assign soundFileAmplitudes [10087] = 8'd113;
   assign soundFileAmplitudes [10088] = 8'd113;
   assign soundFileAmplitudes [10089] = 8'd125;
   assign soundFileAmplitudes [10090] = 8'd131;
   assign soundFileAmplitudes [10091] = 8'd133;
   assign soundFileAmplitudes [10092] = 8'd156;
   assign soundFileAmplitudes [10093] = 8'd167;
   assign soundFileAmplitudes [10094] = 8'd159;
   assign soundFileAmplitudes [10095] = 8'd157;
   assign soundFileAmplitudes [10096] = 8'd151;
   assign soundFileAmplitudes [10097] = 8'd139;
   assign soundFileAmplitudes [10098] = 8'd134;
   assign soundFileAmplitudes [10099] = 8'd136;
   assign soundFileAmplitudes [10100] = 8'd138;
   assign soundFileAmplitudes [10101] = 8'd137;
   assign soundFileAmplitudes [10102] = 8'd125;
   assign soundFileAmplitudes [10103] = 8'd111;
   assign soundFileAmplitudes [10104] = 8'd109;
   assign soundFileAmplitudes [10105] = 8'd116;
   assign soundFileAmplitudes [10106] = 8'd118;
   assign soundFileAmplitudes [10107] = 8'd117;
   assign soundFileAmplitudes [10108] = 8'd113;
   assign soundFileAmplitudes [10109] = 8'd121;
   assign soundFileAmplitudes [10110] = 8'd124;
   assign soundFileAmplitudes [10111] = 8'd107;
   assign soundFileAmplitudes [10112] = 8'd102;
   assign soundFileAmplitudes [10113] = 8'd118;
   assign soundFileAmplitudes [10114] = 8'd122;
   assign soundFileAmplitudes [10115] = 8'd127;
   assign soundFileAmplitudes [10116] = 8'd118;
   assign soundFileAmplitudes [10117] = 8'd112;
   assign soundFileAmplitudes [10118] = 8'd116;
   assign soundFileAmplitudes [10119] = 8'd121;
   assign soundFileAmplitudes [10120] = 8'd133;
   assign soundFileAmplitudes [10121] = 8'd125;
   assign soundFileAmplitudes [10122] = 8'd108;
   assign soundFileAmplitudes [10123] = 8'd110;
   assign soundFileAmplitudes [10124] = 8'd142;
   assign soundFileAmplitudes [10125] = 8'd138;
   assign soundFileAmplitudes [10126] = 8'd134;
   assign soundFileAmplitudes [10127] = 8'd132;
   assign soundFileAmplitudes [10128] = 8'd122;
   assign soundFileAmplitudes [10129] = 8'd118;
   assign soundFileAmplitudes [10130] = 8'd122;
   assign soundFileAmplitudes [10131] = 8'd132;
   assign soundFileAmplitudes [10132] = 8'd145;
   assign soundFileAmplitudes [10133] = 8'd142;
   assign soundFileAmplitudes [10134] = 8'd130;
   assign soundFileAmplitudes [10135] = 8'd129;
   assign soundFileAmplitudes [10136] = 8'd139;
   assign soundFileAmplitudes [10137] = 8'd139;
   assign soundFileAmplitudes [10138] = 8'd134;
   assign soundFileAmplitudes [10139] = 8'd144;
   assign soundFileAmplitudes [10140] = 8'd138;
   assign soundFileAmplitudes [10141] = 8'd135;
   assign soundFileAmplitudes [10142] = 8'd116;
   assign soundFileAmplitudes [10143] = 8'd105;
   assign soundFileAmplitudes [10144] = 8'd113;
   assign soundFileAmplitudes [10145] = 8'd123;
   assign soundFileAmplitudes [10146] = 8'd120;
   assign soundFileAmplitudes [10147] = 8'd109;
   assign soundFileAmplitudes [10148] = 8'd100;
   assign soundFileAmplitudes [10149] = 8'd106;
   assign soundFileAmplitudes [10150] = 8'd113;
   assign soundFileAmplitudes [10151] = 8'd131;
   assign soundFileAmplitudes [10152] = 8'd138;
   assign soundFileAmplitudes [10153] = 8'd134;
   assign soundFileAmplitudes [10154] = 8'd130;
   assign soundFileAmplitudes [10155] = 8'd132;
   assign soundFileAmplitudes [10156] = 8'd148;
   assign soundFileAmplitudes [10157] = 8'd140;
   assign soundFileAmplitudes [10158] = 8'd128;
   assign soundFileAmplitudes [10159] = 8'd114;
   assign soundFileAmplitudes [10160] = 8'd96;
   assign soundFileAmplitudes [10161] = 8'd97;
   assign soundFileAmplitudes [10162] = 8'd103;
   assign soundFileAmplitudes [10163] = 8'd108;
   assign soundFileAmplitudes [10164] = 8'd115;
   assign soundFileAmplitudes [10165] = 8'd107;
   assign soundFileAmplitudes [10166] = 8'd114;
   assign soundFileAmplitudes [10167] = 8'd127;
   assign soundFileAmplitudes [10168] = 8'd156;
   assign soundFileAmplitudes [10169] = 8'd162;
   assign soundFileAmplitudes [10170] = 8'd165;
   assign soundFileAmplitudes [10171] = 8'd160;
   assign soundFileAmplitudes [10172] = 8'd167;
   assign soundFileAmplitudes [10173] = 8'd174;
   assign soundFileAmplitudes [10174] = 8'd157;
   assign soundFileAmplitudes [10175] = 8'd157;
   assign soundFileAmplitudes [10176] = 8'd146;
   assign soundFileAmplitudes [10177] = 8'd138;
   assign soundFileAmplitudes [10178] = 8'd117;
   assign soundFileAmplitudes [10179] = 8'd100;
   assign soundFileAmplitudes [10180] = 8'd86;
   assign soundFileAmplitudes [10181] = 8'd86;
   assign soundFileAmplitudes [10182] = 8'd94;
   assign soundFileAmplitudes [10183] = 8'd105;
   assign soundFileAmplitudes [10184] = 8'd109;
   assign soundFileAmplitudes [10185] = 8'd104;
   assign soundFileAmplitudes [10186] = 8'd106;
   assign soundFileAmplitudes [10187] = 8'd123;
   assign soundFileAmplitudes [10188] = 8'd149;
   assign soundFileAmplitudes [10189] = 8'd155;
   assign soundFileAmplitudes [10190] = 8'd144;
   assign soundFileAmplitudes [10191] = 8'd140;
   assign soundFileAmplitudes [10192] = 8'd127;
   assign soundFileAmplitudes [10193] = 8'd121;
   assign soundFileAmplitudes [10194] = 8'd105;
   assign soundFileAmplitudes [10195] = 8'd88;
   assign soundFileAmplitudes [10196] = 8'd91;
   assign soundFileAmplitudes [10197] = 8'd86;
   assign soundFileAmplitudes [10198] = 8'd102;
   assign soundFileAmplitudes [10199] = 8'd113;
   assign soundFileAmplitudes [10200] = 8'd115;
   assign soundFileAmplitudes [10201] = 8'd116;
   assign soundFileAmplitudes [10202] = 8'd125;
   assign soundFileAmplitudes [10203] = 8'd144;
   assign soundFileAmplitudes [10204] = 8'd179;
   assign soundFileAmplitudes [10205] = 8'd177;
   assign soundFileAmplitudes [10206] = 8'd164;
   assign soundFileAmplitudes [10207] = 8'd169;
   assign soundFileAmplitudes [10208] = 8'd170;
   assign soundFileAmplitudes [10209] = 8'd175;
   assign soundFileAmplitudes [10210] = 8'd162;
   assign soundFileAmplitudes [10211] = 8'd143;
   assign soundFileAmplitudes [10212] = 8'd122;
   assign soundFileAmplitudes [10213] = 8'd113;
   assign soundFileAmplitudes [10214] = 8'd109;
   assign soundFileAmplitudes [10215] = 8'd104;
   assign soundFileAmplitudes [10216] = 8'd107;
   assign soundFileAmplitudes [10217] = 8'd99;
   assign soundFileAmplitudes [10218] = 8'd104;
   assign soundFileAmplitudes [10219] = 8'd111;
   assign soundFileAmplitudes [10220] = 8'd110;
   assign soundFileAmplitudes [10221] = 8'd119;
   assign soundFileAmplitudes [10222] = 8'd119;
   assign soundFileAmplitudes [10223] = 8'd126;
   assign soundFileAmplitudes [10224] = 8'd116;
   assign soundFileAmplitudes [10225] = 8'd109;
   assign soundFileAmplitudes [10226] = 8'd117;
   assign soundFileAmplitudes [10227] = 8'd134;
   assign soundFileAmplitudes [10228] = 8'd137;
   assign soundFileAmplitudes [10229] = 8'd116;
   assign soundFileAmplitudes [10230] = 8'd84;
   assign soundFileAmplitudes [10231] = 8'd92;
   assign soundFileAmplitudes [10232] = 8'd106;
   assign soundFileAmplitudes [10233] = 8'd104;
   assign soundFileAmplitudes [10234] = 8'd117;
   assign soundFileAmplitudes [10235] = 8'd109;
   assign soundFileAmplitudes [10236] = 8'd126;
   assign soundFileAmplitudes [10237] = 8'd128;
   assign soundFileAmplitudes [10238] = 8'd127;
   assign soundFileAmplitudes [10239] = 8'd151;
   assign soundFileAmplitudes [10240] = 8'd177;
   assign soundFileAmplitudes [10241] = 8'd176;
   assign soundFileAmplitudes [10242] = 8'd165;
   assign soundFileAmplitudes [10243] = 8'd161;
   assign soundFileAmplitudes [10244] = 8'd150;
   assign soundFileAmplitudes [10245] = 8'd143;
   assign soundFileAmplitudes [10246] = 8'd141;
   assign soundFileAmplitudes [10247] = 8'd135;
   assign soundFileAmplitudes [10248] = 8'd125;
   assign soundFileAmplitudes [10249] = 8'd115;
   assign soundFileAmplitudes [10250] = 8'd112;
   assign soundFileAmplitudes [10251] = 8'd119;
   assign soundFileAmplitudes [10252] = 8'd120;
   assign soundFileAmplitudes [10253] = 8'd127;
   assign soundFileAmplitudes [10254] = 8'd127;
   assign soundFileAmplitudes [10255] = 8'd123;
   assign soundFileAmplitudes [10256] = 8'd98;
   assign soundFileAmplitudes [10257] = 8'd84;
   assign soundFileAmplitudes [10258] = 8'd103;
   assign soundFileAmplitudes [10259] = 8'd115;
   assign soundFileAmplitudes [10260] = 8'd114;
   assign soundFileAmplitudes [10261] = 8'd111;
   assign soundFileAmplitudes [10262] = 8'd111;
   assign soundFileAmplitudes [10263] = 8'd118;
   assign soundFileAmplitudes [10264] = 8'd109;
   assign soundFileAmplitudes [10265] = 8'd103;
   assign soundFileAmplitudes [10266] = 8'd117;
   assign soundFileAmplitudes [10267] = 8'd127;
   assign soundFileAmplitudes [10268] = 8'd123;
   assign soundFileAmplitudes [10269] = 8'd128;
   assign soundFileAmplitudes [10270] = 8'd138;
   assign soundFileAmplitudes [10271] = 8'd138;
   assign soundFileAmplitudes [10272] = 8'd140;
   assign soundFileAmplitudes [10273] = 8'd140;
   assign soundFileAmplitudes [10274] = 8'd138;
   assign soundFileAmplitudes [10275] = 8'd147;
   assign soundFileAmplitudes [10276] = 8'd145;
   assign soundFileAmplitudes [10277] = 8'd128;
   assign soundFileAmplitudes [10278] = 8'd130;
   assign soundFileAmplitudes [10279] = 8'd127;
   assign soundFileAmplitudes [10280] = 8'd123;
   assign soundFileAmplitudes [10281] = 8'd134;
   assign soundFileAmplitudes [10282] = 8'd129;
   assign soundFileAmplitudes [10283] = 8'd122;
   assign soundFileAmplitudes [10284] = 8'd125;
   assign soundFileAmplitudes [10285] = 8'd129;
   assign soundFileAmplitudes [10286] = 8'd139;
   assign soundFileAmplitudes [10287] = 8'd142;
   assign soundFileAmplitudes [10288] = 8'd138;
   assign soundFileAmplitudes [10289] = 8'd128;
   assign soundFileAmplitudes [10290] = 8'd116;
   assign soundFileAmplitudes [10291] = 8'd117;
   assign soundFileAmplitudes [10292] = 8'd117;
   assign soundFileAmplitudes [10293] = 8'd118;
   assign soundFileAmplitudes [10294] = 8'd119;
   assign soundFileAmplitudes [10295] = 8'd109;
   assign soundFileAmplitudes [10296] = 8'd113;
   assign soundFileAmplitudes [10297] = 8'd120;
   assign soundFileAmplitudes [10298] = 8'd129;
   assign soundFileAmplitudes [10299] = 8'd129;
   assign soundFileAmplitudes [10300] = 8'd116;
   assign soundFileAmplitudes [10301] = 8'd133;
   assign soundFileAmplitudes [10302] = 8'd141;
   assign soundFileAmplitudes [10303] = 8'd136;
   assign soundFileAmplitudes [10304] = 8'd136;
   assign soundFileAmplitudes [10305] = 8'd136;
   assign soundFileAmplitudes [10306] = 8'd139;
   assign soundFileAmplitudes [10307] = 8'd128;
   assign soundFileAmplitudes [10308] = 8'd117;
   assign soundFileAmplitudes [10309] = 8'd100;
   assign soundFileAmplitudes [10310] = 8'd106;
   assign soundFileAmplitudes [10311] = 8'd117;
   assign soundFileAmplitudes [10312] = 8'd121;
   assign soundFileAmplitudes [10313] = 8'd130;
   assign soundFileAmplitudes [10314] = 8'd131;
   assign soundFileAmplitudes [10315] = 8'd123;
   assign soundFileAmplitudes [10316] = 8'd127;
   assign soundFileAmplitudes [10317] = 8'd132;
   assign soundFileAmplitudes [10318] = 8'd132;
   assign soundFileAmplitudes [10319] = 8'd134;
   assign soundFileAmplitudes [10320] = 8'd120;
   assign soundFileAmplitudes [10321] = 8'd111;
   assign soundFileAmplitudes [10322] = 8'd112;
   assign soundFileAmplitudes [10323] = 8'd131;
   assign soundFileAmplitudes [10324] = 8'd138;
   assign soundFileAmplitudes [10325] = 8'd136;
   assign soundFileAmplitudes [10326] = 8'd121;
   assign soundFileAmplitudes [10327] = 8'd108;
   assign soundFileAmplitudes [10328] = 8'd119;
   assign soundFileAmplitudes [10329] = 8'd130;
   assign soundFileAmplitudes [10330] = 8'd135;
   assign soundFileAmplitudes [10331] = 8'd131;
   assign soundFileAmplitudes [10332] = 8'd130;
   assign soundFileAmplitudes [10333] = 8'd137;
   assign soundFileAmplitudes [10334] = 8'd147;
   assign soundFileAmplitudes [10335] = 8'd134;
   assign soundFileAmplitudes [10336] = 8'd136;
   assign soundFileAmplitudes [10337] = 8'd146;
   assign soundFileAmplitudes [10338] = 8'd143;
   assign soundFileAmplitudes [10339] = 8'd132;
   assign soundFileAmplitudes [10340] = 8'd124;
   assign soundFileAmplitudes [10341] = 8'd117;
   assign soundFileAmplitudes [10342] = 8'd115;
   assign soundFileAmplitudes [10343] = 8'd121;
   assign soundFileAmplitudes [10344] = 8'd113;
   assign soundFileAmplitudes [10345] = 8'd119;
   assign soundFileAmplitudes [10346] = 8'd137;
   assign soundFileAmplitudes [10347] = 8'd137;
   assign soundFileAmplitudes [10348] = 8'd127;
   assign soundFileAmplitudes [10349] = 8'd129;
   assign soundFileAmplitudes [10350] = 8'd120;
   assign soundFileAmplitudes [10351] = 8'd127;
   assign soundFileAmplitudes [10352] = 8'd137;
   assign soundFileAmplitudes [10353] = 8'd121;
   assign soundFileAmplitudes [10354] = 8'd110;
   assign soundFileAmplitudes [10355] = 8'd101;
   assign soundFileAmplitudes [10356] = 8'd102;
   assign soundFileAmplitudes [10357] = 8'd115;
   assign soundFileAmplitudes [10358] = 8'd119;
   assign soundFileAmplitudes [10359] = 8'd122;
   assign soundFileAmplitudes [10360] = 8'd128;
   assign soundFileAmplitudes [10361] = 8'd119;
   assign soundFileAmplitudes [10362] = 8'd124;
   assign soundFileAmplitudes [10363] = 8'd124;
   assign soundFileAmplitudes [10364] = 8'd134;
   assign soundFileAmplitudes [10365] = 8'd137;
   assign soundFileAmplitudes [10366] = 8'd132;
   assign soundFileAmplitudes [10367] = 8'd140;
   assign soundFileAmplitudes [10368] = 8'd144;
   assign soundFileAmplitudes [10369] = 8'd143;
   assign soundFileAmplitudes [10370] = 8'd116;
   assign soundFileAmplitudes [10371] = 8'd114;
   assign soundFileAmplitudes [10372] = 8'd113;
   assign soundFileAmplitudes [10373] = 8'd114;
   assign soundFileAmplitudes [10374] = 8'd114;
   assign soundFileAmplitudes [10375] = 8'd113;
   assign soundFileAmplitudes [10376] = 8'd111;
   assign soundFileAmplitudes [10377] = 8'd103;
   assign soundFileAmplitudes [10378] = 8'd115;
   assign soundFileAmplitudes [10379] = 8'd118;
   assign soundFileAmplitudes [10380] = 8'd132;
   assign soundFileAmplitudes [10381] = 8'd148;
   assign soundFileAmplitudes [10382] = 8'd159;
   assign soundFileAmplitudes [10383] = 8'd149;
   assign soundFileAmplitudes [10384] = 8'd152;
   assign soundFileAmplitudes [10385] = 8'd146;
   assign soundFileAmplitudes [10386] = 8'd126;
   assign soundFileAmplitudes [10387] = 8'd125;
   assign soundFileAmplitudes [10388] = 8'd119;
   assign soundFileAmplitudes [10389] = 8'd118;
   assign soundFileAmplitudes [10390] = 8'd109;
   assign soundFileAmplitudes [10391] = 8'd111;
   assign soundFileAmplitudes [10392] = 8'd110;
   assign soundFileAmplitudes [10393] = 8'd109;
   assign soundFileAmplitudes [10394] = 8'd117;
   assign soundFileAmplitudes [10395] = 8'd122;
   assign soundFileAmplitudes [10396] = 8'd128;
   assign soundFileAmplitudes [10397] = 8'd128;
   assign soundFileAmplitudes [10398] = 8'd131;
   assign soundFileAmplitudes [10399] = 8'd138;
   assign soundFileAmplitudes [10400] = 8'd143;
   assign soundFileAmplitudes [10401] = 8'd141;
   assign soundFileAmplitudes [10402] = 8'd144;
   assign soundFileAmplitudes [10403] = 8'd150;
   assign soundFileAmplitudes [10404] = 8'd127;
   assign soundFileAmplitudes [10405] = 8'd116;
   assign soundFileAmplitudes [10406] = 8'd113;
   assign soundFileAmplitudes [10407] = 8'd105;
   assign soundFileAmplitudes [10408] = 8'd96;
   assign soundFileAmplitudes [10409] = 8'd82;
   assign soundFileAmplitudes [10410] = 8'd88;
   assign soundFileAmplitudes [10411] = 8'd104;
   assign soundFileAmplitudes [10412] = 8'd113;
   assign soundFileAmplitudes [10413] = 8'd126;
   assign soundFileAmplitudes [10414] = 8'd135;
   assign soundFileAmplitudes [10415] = 8'd144;
   assign soundFileAmplitudes [10416] = 8'd169;
   assign soundFileAmplitudes [10417] = 8'd176;
   assign soundFileAmplitudes [10418] = 8'd170;
   assign soundFileAmplitudes [10419] = 8'd151;
   assign soundFileAmplitudes [10420] = 8'd148;
   assign soundFileAmplitudes [10421] = 8'd147;
   assign soundFileAmplitudes [10422] = 8'd142;
   assign soundFileAmplitudes [10423] = 8'd130;
   assign soundFileAmplitudes [10424] = 8'd103;
   assign soundFileAmplitudes [10425] = 8'd81;
   assign soundFileAmplitudes [10426] = 8'd74;
   assign soundFileAmplitudes [10427] = 8'd91;
   assign soundFileAmplitudes [10428] = 8'd117;
   assign soundFileAmplitudes [10429] = 8'd120;
   assign soundFileAmplitudes [10430] = 8'd109;
   assign soundFileAmplitudes [10431] = 8'd117;
   assign soundFileAmplitudes [10432] = 8'd128;
   assign soundFileAmplitudes [10433] = 8'd143;
   assign soundFileAmplitudes [10434] = 8'd158;
   assign soundFileAmplitudes [10435] = 8'd169;
   assign soundFileAmplitudes [10436] = 8'd158;
   assign soundFileAmplitudes [10437] = 8'd160;
   assign soundFileAmplitudes [10438] = 8'd134;
   assign soundFileAmplitudes [10439] = 8'd113;
   assign soundFileAmplitudes [10440] = 8'd110;
   assign soundFileAmplitudes [10441] = 8'd94;
   assign soundFileAmplitudes [10442] = 8'd94;
   assign soundFileAmplitudes [10443] = 8'd92;
   assign soundFileAmplitudes [10444] = 8'd94;
   assign soundFileAmplitudes [10445] = 8'd104;
   assign soundFileAmplitudes [10446] = 8'd117;
   assign soundFileAmplitudes [10447] = 8'd114;
   assign soundFileAmplitudes [10448] = 8'd128;
   assign soundFileAmplitudes [10449] = 8'd136;
   assign soundFileAmplitudes [10450] = 8'd152;
   assign soundFileAmplitudes [10451] = 8'd165;
   assign soundFileAmplitudes [10452] = 8'd163;
   assign soundFileAmplitudes [10453] = 8'd154;
   assign soundFileAmplitudes [10454] = 8'd152;
   assign soundFileAmplitudes [10455] = 8'd148;
   assign soundFileAmplitudes [10456] = 8'd140;
   assign soundFileAmplitudes [10457] = 8'd139;
   assign soundFileAmplitudes [10458] = 8'd122;
   assign soundFileAmplitudes [10459] = 8'd113;
   assign soundFileAmplitudes [10460] = 8'd101;
   assign soundFileAmplitudes [10461] = 8'd97;
   assign soundFileAmplitudes [10462] = 8'd104;
   assign soundFileAmplitudes [10463] = 8'd106;
   assign soundFileAmplitudes [10464] = 8'd109;
   assign soundFileAmplitudes [10465] = 8'd116;
   assign soundFileAmplitudes [10466] = 8'd119;
   assign soundFileAmplitudes [10467] = 8'd140;
   assign soundFileAmplitudes [10468] = 8'd153;
   assign soundFileAmplitudes [10469] = 8'd171;
   assign soundFileAmplitudes [10470] = 8'd166;
   assign soundFileAmplitudes [10471] = 8'd149;
   assign soundFileAmplitudes [10472] = 8'd141;
   assign soundFileAmplitudes [10473] = 8'd108;
   assign soundFileAmplitudes [10474] = 8'd98;
   assign soundFileAmplitudes [10475] = 8'd110;
   assign soundFileAmplitudes [10476] = 8'd113;
   assign soundFileAmplitudes [10477] = 8'd105;
   assign soundFileAmplitudes [10478] = 8'd111;
   assign soundFileAmplitudes [10479] = 8'd100;
   assign soundFileAmplitudes [10480] = 8'd109;
   assign soundFileAmplitudes [10481] = 8'd115;
   assign soundFileAmplitudes [10482] = 8'd115;
   assign soundFileAmplitudes [10483] = 8'd138;
   assign soundFileAmplitudes [10484] = 8'd137;
   assign soundFileAmplitudes [10485] = 8'd133;
   assign soundFileAmplitudes [10486] = 8'd134;
   assign soundFileAmplitudes [10487] = 8'd137;
   assign soundFileAmplitudes [10488] = 8'd139;
   assign soundFileAmplitudes [10489] = 8'd142;
   assign soundFileAmplitudes [10490] = 8'd141;
   assign soundFileAmplitudes [10491] = 8'd141;
   assign soundFileAmplitudes [10492] = 8'd126;
   assign soundFileAmplitudes [10493] = 8'd119;
   assign soundFileAmplitudes [10494] = 8'd117;
   assign soundFileAmplitudes [10495] = 8'd116;
   assign soundFileAmplitudes [10496] = 8'd115;
   assign soundFileAmplitudes [10497] = 8'd118;
   assign soundFileAmplitudes [10498] = 8'd118;
   assign soundFileAmplitudes [10499] = 8'd116;
   assign soundFileAmplitudes [10500] = 8'd118;
   assign soundFileAmplitudes [10501] = 8'd124;
   assign soundFileAmplitudes [10502] = 8'd139;
   assign soundFileAmplitudes [10503] = 8'd139;
   assign soundFileAmplitudes [10504] = 8'd150;
   assign soundFileAmplitudes [10505] = 8'd132;
   assign soundFileAmplitudes [10506] = 8'd133;
   assign soundFileAmplitudes [10507] = 8'd132;
   assign soundFileAmplitudes [10508] = 8'd102;
   assign soundFileAmplitudes [10509] = 8'd100;
   assign soundFileAmplitudes [10510] = 8'd98;
   assign soundFileAmplitudes [10511] = 8'd93;
   assign soundFileAmplitudes [10512] = 8'd106;
   assign soundFileAmplitudes [10513] = 8'd115;
   assign soundFileAmplitudes [10514] = 8'd115;
   assign soundFileAmplitudes [10515] = 8'd124;
   assign soundFileAmplitudes [10516] = 8'd122;
   assign soundFileAmplitudes [10517] = 8'd136;
   assign soundFileAmplitudes [10518] = 8'd147;
   assign soundFileAmplitudes [10519] = 8'd151;
   assign soundFileAmplitudes [10520] = 8'd157;
   assign soundFileAmplitudes [10521] = 8'd153;
   assign soundFileAmplitudes [10522] = 8'd144;
   assign soundFileAmplitudes [10523] = 8'd140;
   assign soundFileAmplitudes [10524] = 8'd136;
   assign soundFileAmplitudes [10525] = 8'd130;
   assign soundFileAmplitudes [10526] = 8'd128;
   assign soundFileAmplitudes [10527] = 8'd118;
   assign soundFileAmplitudes [10528] = 8'd110;
   assign soundFileAmplitudes [10529] = 8'd107;
   assign soundFileAmplitudes [10530] = 8'd113;
   assign soundFileAmplitudes [10531] = 8'd118;
   assign soundFileAmplitudes [10532] = 8'd128;
   assign soundFileAmplitudes [10533] = 8'd121;
   assign soundFileAmplitudes [10534] = 8'd115;
   assign soundFileAmplitudes [10535] = 8'd120;
   assign soundFileAmplitudes [10536] = 8'd124;
   assign soundFileAmplitudes [10537] = 8'd137;
   assign soundFileAmplitudes [10538] = 8'd151;
   assign soundFileAmplitudes [10539] = 8'd140;
   assign soundFileAmplitudes [10540] = 8'd132;
   assign soundFileAmplitudes [10541] = 8'd123;
   assign soundFileAmplitudes [10542] = 8'd95;
   assign soundFileAmplitudes [10543] = 8'd96;
   assign soundFileAmplitudes [10544] = 8'd102;
   assign soundFileAmplitudes [10545] = 8'd105;
   assign soundFileAmplitudes [10546] = 8'd101;
   assign soundFileAmplitudes [10547] = 8'd105;
   assign soundFileAmplitudes [10548] = 8'd110;
   assign soundFileAmplitudes [10549] = 8'd125;
   assign soundFileAmplitudes [10550] = 8'd122;
   assign soundFileAmplitudes [10551] = 8'd121;
   assign soundFileAmplitudes [10552] = 8'd138;
   assign soundFileAmplitudes [10553] = 8'd144;
   assign soundFileAmplitudes [10554] = 8'd162;
   assign soundFileAmplitudes [10555] = 8'd169;
   assign soundFileAmplitudes [10556] = 8'd167;
   assign soundFileAmplitudes [10557] = 8'd153;
   assign soundFileAmplitudes [10558] = 8'd145;
   assign soundFileAmplitudes [10559] = 8'd140;
   assign soundFileAmplitudes [10560] = 8'd138;
   assign soundFileAmplitudes [10561] = 8'd128;
   assign soundFileAmplitudes [10562] = 8'd118;
   assign soundFileAmplitudes [10563] = 8'd106;
   assign soundFileAmplitudes [10564] = 8'd107;
   assign soundFileAmplitudes [10565] = 8'd118;
   assign soundFileAmplitudes [10566] = 8'd128;
   assign soundFileAmplitudes [10567] = 8'd138;
   assign soundFileAmplitudes [10568] = 8'd130;
   assign soundFileAmplitudes [10569] = 8'd130;
   assign soundFileAmplitudes [10570] = 8'd113;
   assign soundFileAmplitudes [10571] = 8'd106;
   assign soundFileAmplitudes [10572] = 8'd113;
   assign soundFileAmplitudes [10573] = 8'd113;
   assign soundFileAmplitudes [10574] = 8'd111;
   assign soundFileAmplitudes [10575] = 8'd120;
   assign soundFileAmplitudes [10576] = 8'd124;
   assign soundFileAmplitudes [10577] = 8'd111;
   assign soundFileAmplitudes [10578] = 8'd101;
   assign soundFileAmplitudes [10579] = 8'd106;
   assign soundFileAmplitudes [10580] = 8'd112;
   assign soundFileAmplitudes [10581] = 8'd118;
   assign soundFileAmplitudes [10582] = 8'd121;
   assign soundFileAmplitudes [10583] = 8'd119;
   assign soundFileAmplitudes [10584] = 8'd135;
   assign soundFileAmplitudes [10585] = 8'd131;
   assign soundFileAmplitudes [10586] = 8'd137;
   assign soundFileAmplitudes [10587] = 8'd144;
   assign soundFileAmplitudes [10588] = 8'd152;
   assign soundFileAmplitudes [10589] = 8'd160;
   assign soundFileAmplitudes [10590] = 8'd149;
   assign soundFileAmplitudes [10591] = 8'd149;
   assign soundFileAmplitudes [10592] = 8'd145;
   assign soundFileAmplitudes [10593] = 8'd147;
   assign soundFileAmplitudes [10594] = 8'd148;
   assign soundFileAmplitudes [10595] = 8'd147;
   assign soundFileAmplitudes [10596] = 8'd138;
   assign soundFileAmplitudes [10597] = 8'd133;
   assign soundFileAmplitudes [10598] = 8'd130;
   assign soundFileAmplitudes [10599] = 8'd123;
   assign soundFileAmplitudes [10600] = 8'd127;
   assign soundFileAmplitudes [10601] = 8'd138;
   assign soundFileAmplitudes [10602] = 8'd134;
   assign soundFileAmplitudes [10603] = 8'd128;
   assign soundFileAmplitudes [10604] = 8'd103;
   assign soundFileAmplitudes [10605] = 8'd91;
   assign soundFileAmplitudes [10606] = 8'd86;
   assign soundFileAmplitudes [10607] = 8'd75;
   assign soundFileAmplitudes [10608] = 8'd97;
   assign soundFileAmplitudes [10609] = 8'd108;
   assign soundFileAmplitudes [10610] = 8'd113;
   assign soundFileAmplitudes [10611] = 8'd104;
   assign soundFileAmplitudes [10612] = 8'd90;
   assign soundFileAmplitudes [10613] = 8'd114;
   assign soundFileAmplitudes [10614] = 8'd134;
   assign soundFileAmplitudes [10615] = 8'd138;
   assign soundFileAmplitudes [10616] = 8'd134;
   assign soundFileAmplitudes [10617] = 8'd128;
   assign soundFileAmplitudes [10618] = 8'd136;
   assign soundFileAmplitudes [10619] = 8'd129;
   assign soundFileAmplitudes [10620] = 8'd135;
   assign soundFileAmplitudes [10621] = 8'd136;
   assign soundFileAmplitudes [10622] = 8'd123;
   assign soundFileAmplitudes [10623] = 8'd128;
   assign soundFileAmplitudes [10624] = 8'd136;
   assign soundFileAmplitudes [10625] = 8'd147;
   assign soundFileAmplitudes [10626] = 8'd156;
   assign soundFileAmplitudes [10627] = 8'd154;
   assign soundFileAmplitudes [10628] = 8'd148;
   assign soundFileAmplitudes [10629] = 8'd147;
   assign soundFileAmplitudes [10630] = 8'd142;
   assign soundFileAmplitudes [10631] = 8'd123;
   assign soundFileAmplitudes [10632] = 8'd126;
   assign soundFileAmplitudes [10633] = 8'd131;
   assign soundFileAmplitudes [10634] = 8'd141;
   assign soundFileAmplitudes [10635] = 8'd137;
   assign soundFileAmplitudes [10636] = 8'd107;
   assign soundFileAmplitudes [10637] = 8'd96;
   assign soundFileAmplitudes [10638] = 8'd94;
   assign soundFileAmplitudes [10639] = 8'd101;
   assign soundFileAmplitudes [10640] = 8'd108;
   assign soundFileAmplitudes [10641] = 8'd117;
   assign soundFileAmplitudes [10642] = 8'd120;
   assign soundFileAmplitudes [10643] = 8'd124;
   assign soundFileAmplitudes [10644] = 8'd126;
   assign soundFileAmplitudes [10645] = 8'd126;
   assign soundFileAmplitudes [10646] = 8'd117;
   assign soundFileAmplitudes [10647] = 8'd122;
   assign soundFileAmplitudes [10648] = 8'd119;
   assign soundFileAmplitudes [10649] = 8'd110;
   assign soundFileAmplitudes [10650] = 8'd116;
   assign soundFileAmplitudes [10651] = 8'd109;
   assign soundFileAmplitudes [10652] = 8'd106;
   assign soundFileAmplitudes [10653] = 8'd115;
   assign soundFileAmplitudes [10654] = 8'd130;
   assign soundFileAmplitudes [10655] = 8'd150;
   assign soundFileAmplitudes [10656] = 8'd152;
   assign soundFileAmplitudes [10657] = 8'd143;
   assign soundFileAmplitudes [10658] = 8'd151;
   assign soundFileAmplitudes [10659] = 8'd149;
   assign soundFileAmplitudes [10660] = 8'd156;
   assign soundFileAmplitudes [10661] = 8'd145;
   assign soundFileAmplitudes [10662] = 8'd129;
   assign soundFileAmplitudes [10663] = 8'd120;
   assign soundFileAmplitudes [10664] = 8'd125;
   assign soundFileAmplitudes [10665] = 8'd113;
   assign soundFileAmplitudes [10666] = 8'd106;
   assign soundFileAmplitudes [10667] = 8'd114;
   assign soundFileAmplitudes [10668] = 8'd107;
   assign soundFileAmplitudes [10669] = 8'd107;
   assign soundFileAmplitudes [10670] = 8'd108;
   assign soundFileAmplitudes [10671] = 8'd115;
   assign soundFileAmplitudes [10672] = 8'd123;
   assign soundFileAmplitudes [10673] = 8'd131;
   assign soundFileAmplitudes [10674] = 8'd127;
   assign soundFileAmplitudes [10675] = 8'd136;
   assign soundFileAmplitudes [10676] = 8'd156;
   assign soundFileAmplitudes [10677] = 8'd148;
   assign soundFileAmplitudes [10678] = 8'd137;
   assign soundFileAmplitudes [10679] = 8'd141;
   assign soundFileAmplitudes [10680] = 8'd114;
   assign soundFileAmplitudes [10681] = 8'd93;
   assign soundFileAmplitudes [10682] = 8'd94;
   assign soundFileAmplitudes [10683] = 8'd96;
   assign soundFileAmplitudes [10684] = 8'd104;
   assign soundFileAmplitudes [10685] = 8'd108;
   assign soundFileAmplitudes [10686] = 8'd111;
   assign soundFileAmplitudes [10687] = 8'd128;
   assign soundFileAmplitudes [10688] = 8'd132;
   assign soundFileAmplitudes [10689] = 8'd136;
   assign soundFileAmplitudes [10690] = 8'd148;
   assign soundFileAmplitudes [10691] = 8'd147;
   assign soundFileAmplitudes [10692] = 8'd149;
   assign soundFileAmplitudes [10693] = 8'd157;
   assign soundFileAmplitudes [10694] = 8'd144;
   assign soundFileAmplitudes [10695] = 8'd122;
   assign soundFileAmplitudes [10696] = 8'd120;
   assign soundFileAmplitudes [10697] = 8'd137;
   assign soundFileAmplitudes [10698] = 8'd139;
   assign soundFileAmplitudes [10699] = 8'd118;
   assign soundFileAmplitudes [10700] = 8'd101;
   assign soundFileAmplitudes [10701] = 8'd96;
   assign soundFileAmplitudes [10702] = 8'd116;
   assign soundFileAmplitudes [10703] = 8'd122;
   assign soundFileAmplitudes [10704] = 8'd128;
   assign soundFileAmplitudes [10705] = 8'd133;
   assign soundFileAmplitudes [10706] = 8'd128;
   assign soundFileAmplitudes [10707] = 8'd130;
   assign soundFileAmplitudes [10708] = 8'd134;
   assign soundFileAmplitudes [10709] = 8'd139;
   assign soundFileAmplitudes [10710] = 8'd138;
   assign soundFileAmplitudes [10711] = 8'd130;
   assign soundFileAmplitudes [10712] = 8'd139;
   assign soundFileAmplitudes [10713] = 8'd149;
   assign soundFileAmplitudes [10714] = 8'd141;
   assign soundFileAmplitudes [10715] = 8'd126;
   assign soundFileAmplitudes [10716] = 8'd115;
   assign soundFileAmplitudes [10717] = 8'd116;
   assign soundFileAmplitudes [10718] = 8'd116;
   assign soundFileAmplitudes [10719] = 8'd118;
   assign soundFileAmplitudes [10720] = 8'd117;
   assign soundFileAmplitudes [10721] = 8'd116;
   assign soundFileAmplitudes [10722] = 8'd114;
   assign soundFileAmplitudes [10723] = 8'd108;
   assign soundFileAmplitudes [10724] = 8'd106;
   assign soundFileAmplitudes [10725] = 8'd114;
   assign soundFileAmplitudes [10726] = 8'd121;
   assign soundFileAmplitudes [10727] = 8'd133;
   assign soundFileAmplitudes [10728] = 8'd144;
   assign soundFileAmplitudes [10729] = 8'd144;
   assign soundFileAmplitudes [10730] = 8'd153;
   assign soundFileAmplitudes [10731] = 8'd160;
   assign soundFileAmplitudes [10732] = 8'd133;
   assign soundFileAmplitudes [10733] = 8'd124;
   assign soundFileAmplitudes [10734] = 8'd137;
   assign soundFileAmplitudes [10735] = 8'd133;
   assign soundFileAmplitudes [10736] = 8'd120;
   assign soundFileAmplitudes [10737] = 8'd108;
   assign soundFileAmplitudes [10738] = 8'd116;
   assign soundFileAmplitudes [10739] = 8'd116;
   assign soundFileAmplitudes [10740] = 8'd104;
   assign soundFileAmplitudes [10741] = 8'd103;
   assign soundFileAmplitudes [10742] = 8'd115;
   assign soundFileAmplitudes [10743] = 8'd127;
   assign soundFileAmplitudes [10744] = 8'd124;
   assign soundFileAmplitudes [10745] = 8'd115;
   assign soundFileAmplitudes [10746] = 8'd123;
   assign soundFileAmplitudes [10747] = 8'd141;
   assign soundFileAmplitudes [10748] = 8'd138;
   assign soundFileAmplitudes [10749] = 8'd127;
   assign soundFileAmplitudes [10750] = 8'd126;
   assign soundFileAmplitudes [10751] = 8'd123;
   assign soundFileAmplitudes [10752] = 8'd125;
   assign soundFileAmplitudes [10753] = 8'd108;
   assign soundFileAmplitudes [10754] = 8'd95;
   assign soundFileAmplitudes [10755] = 8'd112;
   assign soundFileAmplitudes [10756] = 8'd125;
   assign soundFileAmplitudes [10757] = 8'd128;
   assign soundFileAmplitudes [10758] = 8'd127;
   assign soundFileAmplitudes [10759] = 8'd132;
   assign soundFileAmplitudes [10760] = 8'd155;
   assign soundFileAmplitudes [10761] = 8'd165;
   assign soundFileAmplitudes [10762] = 8'd174;
   assign soundFileAmplitudes [10763] = 8'd171;
   assign soundFileAmplitudes [10764] = 8'd154;
   assign soundFileAmplitudes [10765] = 8'd143;
   assign soundFileAmplitudes [10766] = 8'd134;
   assign soundFileAmplitudes [10767] = 8'd135;
   assign soundFileAmplitudes [10768] = 8'd115;
   assign soundFileAmplitudes [10769] = 8'd91;
   assign soundFileAmplitudes [10770] = 8'd92;
   assign soundFileAmplitudes [10771] = 8'd112;
   assign soundFileAmplitudes [10772] = 8'd121;
   assign soundFileAmplitudes [10773] = 8'd118;
   assign soundFileAmplitudes [10774] = 8'd120;
   assign soundFileAmplitudes [10775] = 8'd116;
   assign soundFileAmplitudes [10776] = 8'd118;
   assign soundFileAmplitudes [10777] = 8'd109;
   assign soundFileAmplitudes [10778] = 8'd114;
   assign soundFileAmplitudes [10779] = 8'd121;
   assign soundFileAmplitudes [10780] = 8'd116;
   assign soundFileAmplitudes [10781] = 8'd116;
   assign soundFileAmplitudes [10782] = 8'd108;
   assign soundFileAmplitudes [10783] = 8'd112;
   assign soundFileAmplitudes [10784] = 8'd111;
   assign soundFileAmplitudes [10785] = 8'd104;
   assign soundFileAmplitudes [10786] = 8'd109;
   assign soundFileAmplitudes [10787] = 8'd115;
   assign soundFileAmplitudes [10788] = 8'd118;
   assign soundFileAmplitudes [10789] = 8'd128;
   assign soundFileAmplitudes [10790] = 8'd142;
   assign soundFileAmplitudes [10791] = 8'd146;
   assign soundFileAmplitudes [10792] = 8'd157;
   assign soundFileAmplitudes [10793] = 8'd162;
   assign soundFileAmplitudes [10794] = 8'd161;
   assign soundFileAmplitudes [10795] = 8'd148;
   assign soundFileAmplitudes [10796] = 8'd125;
   assign soundFileAmplitudes [10797] = 8'd141;
   assign soundFileAmplitudes [10798] = 8'd142;
   assign soundFileAmplitudes [10799] = 8'd135;
   assign soundFileAmplitudes [10800] = 8'd135;
   assign soundFileAmplitudes [10801] = 8'd134;
   assign soundFileAmplitudes [10802] = 8'd124;
   assign soundFileAmplitudes [10803] = 8'd112;
   assign soundFileAmplitudes [10804] = 8'd105;
   assign soundFileAmplitudes [10805] = 8'd110;
   assign soundFileAmplitudes [10806] = 8'd127;
   assign soundFileAmplitudes [10807] = 8'd118;
   assign soundFileAmplitudes [10808] = 8'd118;
   assign soundFileAmplitudes [10809] = 8'd99;
   assign soundFileAmplitudes [10810] = 8'd98;
   assign soundFileAmplitudes [10811] = 8'd96;
   assign soundFileAmplitudes [10812] = 8'd92;
   assign soundFileAmplitudes [10813] = 8'd107;
   assign soundFileAmplitudes [10814] = 8'd119;
   assign soundFileAmplitudes [10815] = 8'd128;
   assign soundFileAmplitudes [10816] = 8'd114;
   assign soundFileAmplitudes [10817] = 8'd109;
   assign soundFileAmplitudes [10818] = 8'd119;
   assign soundFileAmplitudes [10819] = 8'd142;
   assign soundFileAmplitudes [10820] = 8'd153;
   assign soundFileAmplitudes [10821] = 8'd145;
   assign soundFileAmplitudes [10822] = 8'd148;
   assign soundFileAmplitudes [10823] = 8'd157;
   assign soundFileAmplitudes [10824] = 8'd134;
   assign soundFileAmplitudes [10825] = 8'd133;
   assign soundFileAmplitudes [10826] = 8'd127;
   assign soundFileAmplitudes [10827] = 8'd107;
   assign soundFileAmplitudes [10828] = 8'd104;
   assign soundFileAmplitudes [10829] = 8'd115;
   assign soundFileAmplitudes [10830] = 8'd140;
   assign soundFileAmplitudes [10831] = 8'd141;
   assign soundFileAmplitudes [10832] = 8'd138;
   assign soundFileAmplitudes [10833] = 8'd135;
   assign soundFileAmplitudes [10834] = 8'd150;
   assign soundFileAmplitudes [10835] = 8'd159;
   assign soundFileAmplitudes [10836] = 8'd158;
   assign soundFileAmplitudes [10837] = 8'd163;
   assign soundFileAmplitudes [10838] = 8'd144;
   assign soundFileAmplitudes [10839] = 8'd139;
   assign soundFileAmplitudes [10840] = 8'd102;
   assign soundFileAmplitudes [10841] = 8'd80;
   assign soundFileAmplitudes [10842] = 8'd87;
   assign soundFileAmplitudes [10843] = 8'd98;
   assign soundFileAmplitudes [10844] = 8'd111;
   assign soundFileAmplitudes [10845] = 8'd107;
   assign soundFileAmplitudes [10846] = 8'd118;
   assign soundFileAmplitudes [10847] = 8'd111;
   assign soundFileAmplitudes [10848] = 8'd119;
   assign soundFileAmplitudes [10849] = 8'd116;
   assign soundFileAmplitudes [10850] = 8'd121;
   assign soundFileAmplitudes [10851] = 8'd143;
   assign soundFileAmplitudes [10852] = 8'd153;
   assign soundFileAmplitudes [10853] = 8'd133;
   assign soundFileAmplitudes [10854] = 8'd139;
   assign soundFileAmplitudes [10855] = 8'd150;
   assign soundFileAmplitudes [10856] = 8'd120;
   assign soundFileAmplitudes [10857] = 8'd118;
   assign soundFileAmplitudes [10858] = 8'd107;
   assign soundFileAmplitudes [10859] = 8'd113;
   assign soundFileAmplitudes [10860] = 8'd129;
   assign soundFileAmplitudes [10861] = 8'd123;
   assign soundFileAmplitudes [10862] = 8'd119;
   assign soundFileAmplitudes [10863] = 8'd111;
   assign soundFileAmplitudes [10864] = 8'd108;
   assign soundFileAmplitudes [10865] = 8'd123;
   assign soundFileAmplitudes [10866] = 8'd142;
   assign soundFileAmplitudes [10867] = 8'd145;
   assign soundFileAmplitudes [10868] = 8'd136;
   assign soundFileAmplitudes [10869] = 8'd126;
   assign soundFileAmplitudes [10870] = 8'd115;
   assign soundFileAmplitudes [10871] = 8'd138;
   assign soundFileAmplitudes [10872] = 8'd150;
   assign soundFileAmplitudes [10873] = 8'd148;
   assign soundFileAmplitudes [10874] = 8'd152;
   assign soundFileAmplitudes [10875] = 8'd151;
   assign soundFileAmplitudes [10876] = 8'd156;
   assign soundFileAmplitudes [10877] = 8'd168;
   assign soundFileAmplitudes [10878] = 8'd149;
   assign soundFileAmplitudes [10879] = 8'd119;
   assign soundFileAmplitudes [10880] = 8'd112;
   assign soundFileAmplitudes [10881] = 8'd112;
   assign soundFileAmplitudes [10882] = 8'd111;
   assign soundFileAmplitudes [10883] = 8'd105;
   assign soundFileAmplitudes [10884] = 8'd95;
   assign soundFileAmplitudes [10885] = 8'd80;
   assign soundFileAmplitudes [10886] = 8'd94;
   assign soundFileAmplitudes [10887] = 8'd106;
   assign soundFileAmplitudes [10888] = 8'd124;
   assign soundFileAmplitudes [10889] = 8'd132;
   assign soundFileAmplitudes [10890] = 8'd128;
   assign soundFileAmplitudes [10891] = 8'd130;
   assign soundFileAmplitudes [10892] = 8'd128;
   assign soundFileAmplitudes [10893] = 8'd130;
   assign soundFileAmplitudes [10894] = 8'd125;
   assign soundFileAmplitudes [10895] = 8'd112;
   assign soundFileAmplitudes [10896] = 8'd116;
   assign soundFileAmplitudes [10897] = 8'd124;
   assign soundFileAmplitudes [10898] = 8'd124;
   assign soundFileAmplitudes [10899] = 8'd118;
   assign soundFileAmplitudes [10900] = 8'd89;
   assign soundFileAmplitudes [10901] = 8'd76;
   assign soundFileAmplitudes [10902] = 8'd93;
   assign soundFileAmplitudes [10903] = 8'd135;
   assign soundFileAmplitudes [10904] = 8'd141;
   assign soundFileAmplitudes [10905] = 8'd151;
   assign soundFileAmplitudes [10906] = 8'd157;
   assign soundFileAmplitudes [10907] = 8'd152;
   assign soundFileAmplitudes [10908] = 8'd173;
   assign soundFileAmplitudes [10909] = 8'd170;
   assign soundFileAmplitudes [10910] = 8'd167;
   assign soundFileAmplitudes [10911] = 8'd158;
   assign soundFileAmplitudes [10912] = 8'd139;
   assign soundFileAmplitudes [10913] = 8'd130;
   assign soundFileAmplitudes [10914] = 8'd135;
   assign soundFileAmplitudes [10915] = 8'd130;
   assign soundFileAmplitudes [10916] = 8'd98;
   assign soundFileAmplitudes [10917] = 8'd92;
   assign soundFileAmplitudes [10918] = 8'd100;
   assign soundFileAmplitudes [10919] = 8'd99;
   assign soundFileAmplitudes [10920] = 8'd101;
   assign soundFileAmplitudes [10921] = 8'd102;
   assign soundFileAmplitudes [10922] = 8'd112;
   assign soundFileAmplitudes [10923] = 8'd128;
   assign soundFileAmplitudes [10924] = 8'd133;
   assign soundFileAmplitudes [10925] = 8'd120;
   assign soundFileAmplitudes [10926] = 8'd134;
   assign soundFileAmplitudes [10927] = 8'd131;
   assign soundFileAmplitudes [10928] = 8'd105;
   assign soundFileAmplitudes [10929] = 8'd109;
   assign soundFileAmplitudes [10930] = 8'd112;
   assign soundFileAmplitudes [10931] = 8'd119;
   assign soundFileAmplitudes [10932] = 8'd117;
   assign soundFileAmplitudes [10933] = 8'd114;
   assign soundFileAmplitudes [10934] = 8'd117;
   assign soundFileAmplitudes [10935] = 8'd122;
   assign soundFileAmplitudes [10936] = 8'd130;
   assign soundFileAmplitudes [10937] = 8'd129;
   assign soundFileAmplitudes [10938] = 8'd136;
   assign soundFileAmplitudes [10939] = 8'd155;
   assign soundFileAmplitudes [10940] = 8'd164;
   assign soundFileAmplitudes [10941] = 8'd154;
   assign soundFileAmplitudes [10942] = 8'd145;
   assign soundFileAmplitudes [10943] = 8'd141;
   assign soundFileAmplitudes [10944] = 8'd134;
   assign soundFileAmplitudes [10945] = 8'd134;
   assign soundFileAmplitudes [10946] = 8'd148;
   assign soundFileAmplitudes [10947] = 8'd156;
   assign soundFileAmplitudes [10948] = 8'd153;
   assign soundFileAmplitudes [10949] = 8'd146;
   assign soundFileAmplitudes [10950] = 8'd127;
   assign soundFileAmplitudes [10951] = 8'd113;
   assign soundFileAmplitudes [10952] = 8'd100;
   assign soundFileAmplitudes [10953] = 8'd107;
   assign soundFileAmplitudes [10954] = 8'd119;
   assign soundFileAmplitudes [10955] = 8'd105;
   assign soundFileAmplitudes [10956] = 8'd87;
   assign soundFileAmplitudes [10957] = 8'd85;
   assign soundFileAmplitudes [10958] = 8'd82;
   assign soundFileAmplitudes [10959] = 8'd90;
   assign soundFileAmplitudes [10960] = 8'd102;
   assign soundFileAmplitudes [10961] = 8'd105;
   assign soundFileAmplitudes [10962] = 8'd123;
   assign soundFileAmplitudes [10963] = 8'd115;
   assign soundFileAmplitudes [10964] = 8'd106;
   assign soundFileAmplitudes [10965] = 8'd125;
   assign soundFileAmplitudes [10966] = 8'd131;
   assign soundFileAmplitudes [10967] = 8'd148;
   assign soundFileAmplitudes [10968] = 8'd151;
   assign soundFileAmplitudes [10969] = 8'd147;
   assign soundFileAmplitudes [10970] = 8'd148;
   assign soundFileAmplitudes [10971] = 8'd140;
   assign soundFileAmplitudes [10972] = 8'd127;
   assign soundFileAmplitudes [10973] = 8'd93;
   assign soundFileAmplitudes [10974] = 8'd110;
   assign soundFileAmplitudes [10975] = 8'd134;
   assign soundFileAmplitudes [10976] = 8'd129;
   assign soundFileAmplitudes [10977] = 8'd151;
   assign soundFileAmplitudes [10978] = 8'd154;
   assign soundFileAmplitudes [10979] = 8'd141;
   assign soundFileAmplitudes [10980] = 8'd140;
   assign soundFileAmplitudes [10981] = 8'd128;
   assign soundFileAmplitudes [10982] = 8'd137;
   assign soundFileAmplitudes [10983] = 8'd153;
   assign soundFileAmplitudes [10984] = 8'd151;
   assign soundFileAmplitudes [10985] = 8'd161;
   assign soundFileAmplitudes [10986] = 8'd162;
   assign soundFileAmplitudes [10987] = 8'd151;
   assign soundFileAmplitudes [10988] = 8'd142;
   assign soundFileAmplitudes [10989] = 8'd125;
   assign soundFileAmplitudes [10990] = 8'd101;
   assign soundFileAmplitudes [10991] = 8'd89;
   assign soundFileAmplitudes [10992] = 8'd82;
   assign soundFileAmplitudes [10993] = 8'd93;
   assign soundFileAmplitudes [10994] = 8'd91;
   assign soundFileAmplitudes [10995] = 8'd86;
   assign soundFileAmplitudes [10996] = 8'd94;
   assign soundFileAmplitudes [10997] = 8'd102;
   assign soundFileAmplitudes [10998] = 8'd104;
   assign soundFileAmplitudes [10999] = 8'd126;
   assign soundFileAmplitudes [11000] = 8'd137;
   assign soundFileAmplitudes [11001] = 8'd127;
   assign soundFileAmplitudes [11002] = 8'd133;
   assign soundFileAmplitudes [11003] = 8'd124;
   assign soundFileAmplitudes [11004] = 8'd129;
   assign soundFileAmplitudes [11005] = 8'd136;
   assign soundFileAmplitudes [11006] = 8'd127;
   assign soundFileAmplitudes [11007] = 8'd99;
   assign soundFileAmplitudes [11008] = 8'd142;
   assign soundFileAmplitudes [11009] = 8'd166;
   assign soundFileAmplitudes [11010] = 8'd146;
   assign soundFileAmplitudes [11011] = 8'd158;
   assign soundFileAmplitudes [11012] = 8'd145;
   assign soundFileAmplitudes [11013] = 8'd133;
   assign soundFileAmplitudes [11014] = 8'd144;
   assign soundFileAmplitudes [11015] = 8'd140;
   assign soundFileAmplitudes [11016] = 8'd133;
   assign soundFileAmplitudes [11017] = 8'd134;
   assign soundFileAmplitudes [11018] = 8'd134;
   assign soundFileAmplitudes [11019] = 8'd144;
   assign soundFileAmplitudes [11020] = 8'd133;
   assign soundFileAmplitudes [11021] = 8'd126;
   assign soundFileAmplitudes [11022] = 8'd107;
   assign soundFileAmplitudes [11023] = 8'd116;
   assign soundFileAmplitudes [11024] = 8'd136;
   assign soundFileAmplitudes [11025] = 8'd132;
   assign soundFileAmplitudes [11026] = 8'd127;
   assign soundFileAmplitudes [11027] = 8'd128;
   assign soundFileAmplitudes [11028] = 8'd115;
   assign soundFileAmplitudes [11029] = 8'd108;
   assign soundFileAmplitudes [11030] = 8'd112;
   assign soundFileAmplitudes [11031] = 8'd116;
   assign soundFileAmplitudes [11032] = 8'd102;
   assign soundFileAmplitudes [11033] = 8'd90;
   assign soundFileAmplitudes [11034] = 8'd92;
   assign soundFileAmplitudes [11035] = 8'd83;
   assign soundFileAmplitudes [11036] = 8'd77;
   assign soundFileAmplitudes [11037] = 8'd83;
   assign soundFileAmplitudes [11038] = 8'd93;
   assign soundFileAmplitudes [11039] = 8'd105;
   assign soundFileAmplitudes [11040] = 8'd116;
   assign soundFileAmplitudes [11041] = 8'd98;
   assign soundFileAmplitudes [11042] = 8'd147;
   assign soundFileAmplitudes [11043] = 8'd179;
   assign soundFileAmplitudes [11044] = 8'd167;
   assign soundFileAmplitudes [11045] = 8'd186;
   assign soundFileAmplitudes [11046] = 8'd185;
   assign soundFileAmplitudes [11047] = 8'd182;
   assign soundFileAmplitudes [11048] = 8'd178;
   assign soundFileAmplitudes [11049] = 8'd171;
   assign soundFileAmplitudes [11050] = 8'd156;
   assign soundFileAmplitudes [11051] = 8'd126;
   assign soundFileAmplitudes [11052] = 8'd119;
   assign soundFileAmplitudes [11053] = 8'd118;
   assign soundFileAmplitudes [11054] = 8'd109;
   assign soundFileAmplitudes [11055] = 8'd114;
   assign soundFileAmplitudes [11056] = 8'd117;
   assign soundFileAmplitudes [11057] = 8'd122;
   assign soundFileAmplitudes [11058] = 8'd118;
   assign soundFileAmplitudes [11059] = 8'd110;
   assign soundFileAmplitudes [11060] = 8'd118;
   assign soundFileAmplitudes [11061] = 8'd123;
   assign soundFileAmplitudes [11062] = 8'd117;
   assign soundFileAmplitudes [11063] = 8'd121;
   assign soundFileAmplitudes [11064] = 8'd123;
   assign soundFileAmplitudes [11065] = 8'd119;
   assign soundFileAmplitudes [11066] = 8'd114;
   assign soundFileAmplitudes [11067] = 8'd113;
   assign soundFileAmplitudes [11068] = 8'd99;
   assign soundFileAmplitudes [11069] = 8'd90;
   assign soundFileAmplitudes [11070] = 8'd91;
   assign soundFileAmplitudes [11071] = 8'd95;
   assign soundFileAmplitudes [11072] = 8'd101;
   assign soundFileAmplitudes [11073] = 8'd94;
   assign soundFileAmplitudes [11074] = 8'd106;
   assign soundFileAmplitudes [11075] = 8'd103;
   assign soundFileAmplitudes [11076] = 8'd116;
   assign soundFileAmplitudes [11077] = 8'd133;
   assign soundFileAmplitudes [11078] = 8'd144;
   assign soundFileAmplitudes [11079] = 8'd154;
   assign soundFileAmplitudes [11080] = 8'd155;
   assign soundFileAmplitudes [11081] = 8'd176;
   assign soundFileAmplitudes [11082] = 8'd177;
   assign soundFileAmplitudes [11083] = 8'd162;
   assign soundFileAmplitudes [11084] = 8'd153;
   assign soundFileAmplitudes [11085] = 8'd151;
   assign soundFileAmplitudes [11086] = 8'd150;
   assign soundFileAmplitudes [11087] = 8'd148;
   assign soundFileAmplitudes [11088] = 8'd146;
   assign soundFileAmplitudes [11089] = 8'd131;
   assign soundFileAmplitudes [11090] = 8'd124;
   assign soundFileAmplitudes [11091] = 8'd115;
   assign soundFileAmplitudes [11092] = 8'd102;
   assign soundFileAmplitudes [11093] = 8'd107;
   assign soundFileAmplitudes [11094] = 8'd109;
   assign soundFileAmplitudes [11095] = 8'd99;
   assign soundFileAmplitudes [11096] = 8'd88;
   assign soundFileAmplitudes [11097] = 8'd103;
   assign soundFileAmplitudes [11098] = 8'd120;
   assign soundFileAmplitudes [11099] = 8'd125;
   assign soundFileAmplitudes [11100] = 8'd132;
   assign soundFileAmplitudes [11101] = 8'd132;
   assign soundFileAmplitudes [11102] = 8'd133;
   assign soundFileAmplitudes [11103] = 8'd127;
   assign soundFileAmplitudes [11104] = 8'd125;
   assign soundFileAmplitudes [11105] = 8'd123;
   assign soundFileAmplitudes [11106] = 8'd116;
   assign soundFileAmplitudes [11107] = 8'd112;
   assign soundFileAmplitudes [11108] = 8'd102;
   assign soundFileAmplitudes [11109] = 8'd88;
   assign soundFileAmplitudes [11110] = 8'd80;
   assign soundFileAmplitudes [11111] = 8'd95;
   assign soundFileAmplitudes [11112] = 8'd117;
   assign soundFileAmplitudes [11113] = 8'd127;
   assign soundFileAmplitudes [11114] = 8'd136;
   assign soundFileAmplitudes [11115] = 8'd149;
   assign soundFileAmplitudes [11116] = 8'd161;
   assign soundFileAmplitudes [11117] = 8'd169;
   assign soundFileAmplitudes [11118] = 8'd178;
   assign soundFileAmplitudes [11119] = 8'd188;
   assign soundFileAmplitudes [11120] = 8'd192;
   assign soundFileAmplitudes [11121] = 8'd168;
   assign soundFileAmplitudes [11122] = 8'd146;
   assign soundFileAmplitudes [11123] = 8'd136;
   assign soundFileAmplitudes [11124] = 8'd133;
   assign soundFileAmplitudes [11125] = 8'd110;
   assign soundFileAmplitudes [11126] = 8'd88;
   assign soundFileAmplitudes [11127] = 8'd96;
   assign soundFileAmplitudes [11128] = 8'd97;
   assign soundFileAmplitudes [11129] = 8'd110;
   assign soundFileAmplitudes [11130] = 8'd105;
   assign soundFileAmplitudes [11131] = 8'd95;
   assign soundFileAmplitudes [11132] = 8'd99;
   assign soundFileAmplitudes [11133] = 8'd102;
   assign soundFileAmplitudes [11134] = 8'd127;
   assign soundFileAmplitudes [11135] = 8'd136;
   assign soundFileAmplitudes [11136] = 8'd128;
   assign soundFileAmplitudes [11137] = 8'd130;
   assign soundFileAmplitudes [11138] = 8'd100;
   assign soundFileAmplitudes [11139] = 8'd83;
   assign soundFileAmplitudes [11140] = 8'd104;
   assign soundFileAmplitudes [11141] = 8'd104;
   assign soundFileAmplitudes [11142] = 8'd108;
   assign soundFileAmplitudes [11143] = 8'd114;
   assign soundFileAmplitudes [11144] = 8'd115;
   assign soundFileAmplitudes [11145] = 8'd128;
   assign soundFileAmplitudes [11146] = 8'd148;
   assign soundFileAmplitudes [11147] = 8'd156;
   assign soundFileAmplitudes [11148] = 8'd152;
   assign soundFileAmplitudes [11149] = 8'd167;
   assign soundFileAmplitudes [11150] = 8'd172;
   assign soundFileAmplitudes [11151] = 8'd167;
   assign soundFileAmplitudes [11152] = 8'd164;
   assign soundFileAmplitudes [11153] = 8'd161;
   assign soundFileAmplitudes [11154] = 8'd143;
   assign soundFileAmplitudes [11155] = 8'd131;
   assign soundFileAmplitudes [11156] = 8'd132;
   assign soundFileAmplitudes [11157] = 8'd136;
   assign soundFileAmplitudes [11158] = 8'd132;
   assign soundFileAmplitudes [11159] = 8'd116;
   assign soundFileAmplitudes [11160] = 8'd114;
   assign soundFileAmplitudes [11161] = 8'd114;
   assign soundFileAmplitudes [11162] = 8'd123;
   assign soundFileAmplitudes [11163] = 8'd127;
   assign soundFileAmplitudes [11164] = 8'd131;
   assign soundFileAmplitudes [11165] = 8'd115;
   assign soundFileAmplitudes [11166] = 8'd98;
   assign soundFileAmplitudes [11167] = 8'd77;
   assign soundFileAmplitudes [11168] = 8'd63;
   assign soundFileAmplitudes [11169] = 8'd82;
   assign soundFileAmplitudes [11170] = 8'd90;
   assign soundFileAmplitudes [11171] = 8'd99;
   assign soundFileAmplitudes [11172] = 8'd113;
   assign soundFileAmplitudes [11173] = 8'd107;
   assign soundFileAmplitudes [11174] = 8'd107;
   assign soundFileAmplitudes [11175] = 8'd129;
   assign soundFileAmplitudes [11176] = 8'd134;
   assign soundFileAmplitudes [11177] = 8'd133;
   assign soundFileAmplitudes [11178] = 8'd143;
   assign soundFileAmplitudes [11179] = 8'd148;
   assign soundFileAmplitudes [11180] = 8'd139;
   assign soundFileAmplitudes [11181] = 8'd131;
   assign soundFileAmplitudes [11182] = 8'd137;
   assign soundFileAmplitudes [11183] = 8'd138;
   assign soundFileAmplitudes [11184] = 8'd124;
   assign soundFileAmplitudes [11185] = 8'd136;
   assign soundFileAmplitudes [11186] = 8'd156;
   assign soundFileAmplitudes [11187] = 8'd168;
   assign soundFileAmplitudes [11188] = 8'd167;
   assign soundFileAmplitudes [11189] = 8'd162;
   assign soundFileAmplitudes [11190] = 8'd149;
   assign soundFileAmplitudes [11191] = 8'd144;
   assign soundFileAmplitudes [11192] = 8'd137;
   assign soundFileAmplitudes [11193] = 8'd139;
   assign soundFileAmplitudes [11194] = 8'd128;
   assign soundFileAmplitudes [11195] = 8'd111;
   assign soundFileAmplitudes [11196] = 8'd106;
   assign soundFileAmplitudes [11197] = 8'd86;
   assign soundFileAmplitudes [11198] = 8'd97;
   assign soundFileAmplitudes [11199] = 8'd93;
   assign soundFileAmplitudes [11200] = 8'd89;
   assign soundFileAmplitudes [11201] = 8'd90;
   assign soundFileAmplitudes [11202] = 8'd87;
   assign soundFileAmplitudes [11203] = 8'd99;
   assign soundFileAmplitudes [11204] = 8'd123;
   assign soundFileAmplitudes [11205] = 8'd124;
   assign soundFileAmplitudes [11206] = 8'd127;
   assign soundFileAmplitudes [11207] = 8'd139;
   assign soundFileAmplitudes [11208] = 8'd131;
   assign soundFileAmplitudes [11209] = 8'd121;
   assign soundFileAmplitudes [11210] = 8'd112;
   assign soundFileAmplitudes [11211] = 8'd130;
   assign soundFileAmplitudes [11212] = 8'd144;
   assign soundFileAmplitudes [11213] = 8'd131;
   assign soundFileAmplitudes [11214] = 8'd113;
   assign soundFileAmplitudes [11215] = 8'd109;
   assign soundFileAmplitudes [11216] = 8'd140;
   assign soundFileAmplitudes [11217] = 8'd154;
   assign soundFileAmplitudes [11218] = 8'd157;
   assign soundFileAmplitudes [11219] = 8'd165;
   assign soundFileAmplitudes [11220] = 8'd161;
   assign soundFileAmplitudes [11221] = 8'd168;
   assign soundFileAmplitudes [11222] = 8'd162;
   assign soundFileAmplitudes [11223] = 8'd169;
   assign soundFileAmplitudes [11224] = 8'd148;
   assign soundFileAmplitudes [11225] = 8'd135;
   assign soundFileAmplitudes [11226] = 8'd109;
   assign soundFileAmplitudes [11227] = 8'd90;
   assign soundFileAmplitudes [11228] = 8'd105;
   assign soundFileAmplitudes [11229] = 8'd102;
   assign soundFileAmplitudes [11230] = 8'd108;
   assign soundFileAmplitudes [11231] = 8'd94;
   assign soundFileAmplitudes [11232] = 8'd84;
   assign soundFileAmplitudes [11233] = 8'd91;
   assign soundFileAmplitudes [11234] = 8'd108;
   assign soundFileAmplitudes [11235] = 8'd129;
   assign soundFileAmplitudes [11236] = 8'd131;
   assign soundFileAmplitudes [11237] = 8'd113;
   assign soundFileAmplitudes [11238] = 8'd125;
   assign soundFileAmplitudes [11239] = 8'd131;
   assign soundFileAmplitudes [11240] = 8'd141;
   assign soundFileAmplitudes [11241] = 8'd142;
   assign soundFileAmplitudes [11242] = 8'd117;
   assign soundFileAmplitudes [11243] = 8'd99;
   assign soundFileAmplitudes [11244] = 8'd91;
   assign soundFileAmplitudes [11245] = 8'd109;
   assign soundFileAmplitudes [11246] = 8'd116;
   assign soundFileAmplitudes [11247] = 8'd96;
   assign soundFileAmplitudes [11248] = 8'd91;
   assign soundFileAmplitudes [11249] = 8'd104;
   assign soundFileAmplitudes [11250] = 8'd126;
   assign soundFileAmplitudes [11251] = 8'd151;
   assign soundFileAmplitudes [11252] = 8'd153;
   assign soundFileAmplitudes [11253] = 8'd170;
   assign soundFileAmplitudes [11254] = 8'd166;
   assign soundFileAmplitudes [11255] = 8'd157;
   assign soundFileAmplitudes [11256] = 8'd145;
   assign soundFileAmplitudes [11257] = 8'd143;
   assign soundFileAmplitudes [11258] = 8'd152;
   assign soundFileAmplitudes [11259] = 8'd142;
   assign soundFileAmplitudes [11260] = 8'd146;
   assign soundFileAmplitudes [11261] = 8'd134;
   assign soundFileAmplitudes [11262] = 8'd125;
   assign soundFileAmplitudes [11263] = 8'd119;
   assign soundFileAmplitudes [11264] = 8'd123;
   assign soundFileAmplitudes [11265] = 8'd142;
   assign soundFileAmplitudes [11266] = 8'd150;
   assign soundFileAmplitudes [11267] = 8'd150;
   assign soundFileAmplitudes [11268] = 8'd143;
   assign soundFileAmplitudes [11269] = 8'd113;
   assign soundFileAmplitudes [11270] = 8'd104;
   assign soundFileAmplitudes [11271] = 8'd110;
   assign soundFileAmplitudes [11272] = 8'd109;
   assign soundFileAmplitudes [11273] = 8'd106;
   assign soundFileAmplitudes [11274] = 8'd105;
   assign soundFileAmplitudes [11275] = 8'd119;
   assign soundFileAmplitudes [11276] = 8'd127;
   assign soundFileAmplitudes [11277] = 8'd132;
   assign soundFileAmplitudes [11278] = 8'd125;
   assign soundFileAmplitudes [11279] = 8'd115;
   assign soundFileAmplitudes [11280] = 8'd102;
   assign soundFileAmplitudes [11281] = 8'd97;
   assign soundFileAmplitudes [11282] = 8'd85;
   assign soundFileAmplitudes [11283] = 8'd100;
   assign soundFileAmplitudes [11284] = 8'd114;
   assign soundFileAmplitudes [11285] = 8'd110;
   assign soundFileAmplitudes [11286] = 8'd95;
   assign soundFileAmplitudes [11287] = 8'd72;
   assign soundFileAmplitudes [11288] = 8'd95;
   assign soundFileAmplitudes [11289] = 8'd120;
   assign soundFileAmplitudes [11290] = 8'd141;
   assign soundFileAmplitudes [11291] = 8'd142;
   assign soundFileAmplitudes [11292] = 8'd153;
   assign soundFileAmplitudes [11293] = 8'd169;
   assign soundFileAmplitudes [11294] = 8'd184;
   assign soundFileAmplitudes [11295] = 8'd188;
   assign soundFileAmplitudes [11296] = 8'd196;
   assign soundFileAmplitudes [11297] = 8'd195;
   assign soundFileAmplitudes [11298] = 8'd180;
   assign soundFileAmplitudes [11299] = 8'd157;
   assign soundFileAmplitudes [11300] = 8'd145;
   assign soundFileAmplitudes [11301] = 8'd141;
   assign soundFileAmplitudes [11302] = 8'd125;
   assign soundFileAmplitudes [11303] = 8'd111;
   assign soundFileAmplitudes [11304] = 8'd90;
   assign soundFileAmplitudes [11305] = 8'd97;
   assign soundFileAmplitudes [11306] = 8'd103;
   assign soundFileAmplitudes [11307] = 8'd106;
   assign soundFileAmplitudes [11308] = 8'd94;
   assign soundFileAmplitudes [11309] = 8'd88;
   assign soundFileAmplitudes [11310] = 8'd96;
   assign soundFileAmplitudes [11311] = 8'd120;
   assign soundFileAmplitudes [11312] = 8'd119;
   assign soundFileAmplitudes [11313] = 8'd121;
   assign soundFileAmplitudes [11314] = 8'd125;
   assign soundFileAmplitudes [11315] = 8'd109;
   assign soundFileAmplitudes [11316] = 8'd100;
   assign soundFileAmplitudes [11317] = 8'd71;
   assign soundFileAmplitudes [11318] = 8'd73;
   assign soundFileAmplitudes [11319] = 8'd85;
   assign soundFileAmplitudes [11320] = 8'd97;
   assign soundFileAmplitudes [11321] = 8'd99;
   assign soundFileAmplitudes [11322] = 8'd109;
   assign soundFileAmplitudes [11323] = 8'd118;
   assign soundFileAmplitudes [11324] = 8'd131;
   assign soundFileAmplitudes [11325] = 8'd150;
   assign soundFileAmplitudes [11326] = 8'd157;
   assign soundFileAmplitudes [11327] = 8'd163;
   assign soundFileAmplitudes [11328] = 8'd180;
   assign soundFileAmplitudes [11329] = 8'd190;
   assign soundFileAmplitudes [11330] = 8'd181;
   assign soundFileAmplitudes [11331] = 8'd188;
   assign soundFileAmplitudes [11332] = 8'd173;
   assign soundFileAmplitudes [11333] = 8'd151;
   assign soundFileAmplitudes [11334] = 8'd135;
   assign soundFileAmplitudes [11335] = 8'd143;
   assign soundFileAmplitudes [11336] = 8'd162;
   assign soundFileAmplitudes [11337] = 8'd152;
   assign soundFileAmplitudes [11338] = 8'd122;
   assign soundFileAmplitudes [11339] = 8'd100;
   assign soundFileAmplitudes [11340] = 8'd96;
   assign soundFileAmplitudes [11341] = 8'd105;
   assign soundFileAmplitudes [11342] = 8'd96;
   assign soundFileAmplitudes [11343] = 8'd87;
   assign soundFileAmplitudes [11344] = 8'd105;
   assign soundFileAmplitudes [11345] = 8'd107;
   assign soundFileAmplitudes [11346] = 8'd102;
   assign soundFileAmplitudes [11347] = 8'd82;
   assign soundFileAmplitudes [11348] = 8'd76;
   assign soundFileAmplitudes [11349] = 8'd94;
   assign soundFileAmplitudes [11350] = 8'd105;
   assign soundFileAmplitudes [11351] = 8'd104;
   assign soundFileAmplitudes [11352] = 8'd93;
   assign soundFileAmplitudes [11353] = 8'd90;
   assign soundFileAmplitudes [11354] = 8'd98;
   assign soundFileAmplitudes [11355] = 8'd107;
   assign soundFileAmplitudes [11356] = 8'd120;
   assign soundFileAmplitudes [11357] = 8'd134;
   assign soundFileAmplitudes [11358] = 8'd147;
   assign soundFileAmplitudes [11359] = 8'd158;
   assign soundFileAmplitudes [11360] = 8'd142;
   assign soundFileAmplitudes [11361] = 8'd139;
   assign soundFileAmplitudes [11362] = 8'd158;
   assign soundFileAmplitudes [11363] = 8'd161;
   assign soundFileAmplitudes [11364] = 8'd157;
   assign soundFileAmplitudes [11365] = 8'd147;
   assign soundFileAmplitudes [11366] = 8'd148;
   assign soundFileAmplitudes [11367] = 8'd177;
   assign soundFileAmplitudes [11368] = 8'd186;
   assign soundFileAmplitudes [11369] = 8'd174;
   assign soundFileAmplitudes [11370] = 8'd158;
   assign soundFileAmplitudes [11371] = 8'd151;
   assign soundFileAmplitudes [11372] = 8'd156;
   assign soundFileAmplitudes [11373] = 8'd144;
   assign soundFileAmplitudes [11374] = 8'd139;
   assign soundFileAmplitudes [11375] = 8'd121;
   assign soundFileAmplitudes [11376] = 8'd101;
   assign soundFileAmplitudes [11377] = 8'd86;
   assign soundFileAmplitudes [11378] = 8'd60;
   assign soundFileAmplitudes [11379] = 8'd64;
   assign soundFileAmplitudes [11380] = 8'd65;
   assign soundFileAmplitudes [11381] = 8'd73;
   assign soundFileAmplitudes [11382] = 8'd90;
   assign soundFileAmplitudes [11383] = 8'd99;
   assign soundFileAmplitudes [11384] = 8'd119;
   assign soundFileAmplitudes [11385] = 8'd128;
   assign soundFileAmplitudes [11386] = 8'd123;
   assign soundFileAmplitudes [11387] = 8'd127;
   assign soundFileAmplitudes [11388] = 8'd139;
   assign soundFileAmplitudes [11389] = 8'd142;
   assign soundFileAmplitudes [11390] = 8'd136;
   assign soundFileAmplitudes [11391] = 8'd125;
   assign soundFileAmplitudes [11392] = 8'd116;
   assign soundFileAmplitudes [11393] = 8'd116;
   assign soundFileAmplitudes [11394] = 8'd121;
   assign soundFileAmplitudes [11395] = 8'd117;
   assign soundFileAmplitudes [11396] = 8'd127;
   assign soundFileAmplitudes [11397] = 8'd133;
   assign soundFileAmplitudes [11398] = 8'd130;
   assign soundFileAmplitudes [11399] = 8'd138;
   assign soundFileAmplitudes [11400] = 8'd151;
   assign soundFileAmplitudes [11401] = 8'd154;
   assign soundFileAmplitudes [11402] = 8'd153;
   assign soundFileAmplitudes [11403] = 8'd141;
   assign soundFileAmplitudes [11404] = 8'd140;
   assign soundFileAmplitudes [11405] = 8'd162;
   assign soundFileAmplitudes [11406] = 8'd164;
   assign soundFileAmplitudes [11407] = 8'd166;
   assign soundFileAmplitudes [11408] = 8'd147;
   assign soundFileAmplitudes [11409] = 8'd120;
   assign soundFileAmplitudes [11410] = 8'd112;
   assign soundFileAmplitudes [11411] = 8'd107;
   assign soundFileAmplitudes [11412] = 8'd104;
   assign soundFileAmplitudes [11413] = 8'd85;
   assign soundFileAmplitudes [11414] = 8'd76;
   assign soundFileAmplitudes [11415] = 8'd92;
   assign soundFileAmplitudes [11416] = 8'd101;
   assign soundFileAmplitudes [11417] = 8'd112;
   assign soundFileAmplitudes [11418] = 8'd124;
   assign soundFileAmplitudes [11419] = 8'd127;
   assign soundFileAmplitudes [11420] = 8'd144;
   assign soundFileAmplitudes [11421] = 8'd152;
   assign soundFileAmplitudes [11422] = 8'd139;
   assign soundFileAmplitudes [11423] = 8'd126;
   assign soundFileAmplitudes [11424] = 8'd125;
   assign soundFileAmplitudes [11425] = 8'd112;
   assign soundFileAmplitudes [11426] = 8'd86;
   assign soundFileAmplitudes [11427] = 8'd96;
   assign soundFileAmplitudes [11428] = 8'd116;
   assign soundFileAmplitudes [11429] = 8'd124;
   assign soundFileAmplitudes [11430] = 8'd124;
   assign soundFileAmplitudes [11431] = 8'd117;
   assign soundFileAmplitudes [11432] = 8'd117;
   assign soundFileAmplitudes [11433] = 8'd129;
   assign soundFileAmplitudes [11434] = 8'd141;
   assign soundFileAmplitudes [11435] = 8'd139;
   assign soundFileAmplitudes [11436] = 8'd145;
   assign soundFileAmplitudes [11437] = 8'd154;
   assign soundFileAmplitudes [11438] = 8'd157;
   assign soundFileAmplitudes [11439] = 8'd145;
   assign soundFileAmplitudes [11440] = 8'd129;
   assign soundFileAmplitudes [11441] = 8'd132;
   assign soundFileAmplitudes [11442] = 8'd131;
   assign soundFileAmplitudes [11443] = 8'd143;
   assign soundFileAmplitudes [11444] = 8'd152;
   assign soundFileAmplitudes [11445] = 8'd133;
   assign soundFileAmplitudes [11446] = 8'd123;
   assign soundFileAmplitudes [11447] = 8'd112;
   assign soundFileAmplitudes [11448] = 8'd115;
   assign soundFileAmplitudes [11449] = 8'd130;
   assign soundFileAmplitudes [11450] = 8'd133;
   assign soundFileAmplitudes [11451] = 8'd131;
   assign soundFileAmplitudes [11452] = 8'd132;
   assign soundFileAmplitudes [11453] = 8'd130;
   assign soundFileAmplitudes [11454] = 8'd123;
   assign soundFileAmplitudes [11455] = 8'd120;
   assign soundFileAmplitudes [11456] = 8'd119;
   assign soundFileAmplitudes [11457] = 8'd111;
   assign soundFileAmplitudes [11458] = 8'd101;
   assign soundFileAmplitudes [11459] = 8'd106;
   assign soundFileAmplitudes [11460] = 8'd111;
   assign soundFileAmplitudes [11461] = 8'd118;
   assign soundFileAmplitudes [11462] = 8'd110;
   assign soundFileAmplitudes [11463] = 8'd103;
   assign soundFileAmplitudes [11464] = 8'd112;
   assign soundFileAmplitudes [11465] = 8'd114;
   assign soundFileAmplitudes [11466] = 8'd119;
   assign soundFileAmplitudes [11467] = 8'd138;
   assign soundFileAmplitudes [11468] = 8'd146;
   assign soundFileAmplitudes [11469] = 8'd143;
   assign soundFileAmplitudes [11470] = 8'd134;
   assign soundFileAmplitudes [11471] = 8'd113;
   assign soundFileAmplitudes [11472] = 8'd109;
   assign soundFileAmplitudes [11473] = 8'd119;
   assign soundFileAmplitudes [11474] = 8'd132;
   assign soundFileAmplitudes [11475] = 8'd125;
   assign soundFileAmplitudes [11476] = 8'd124;
   assign soundFileAmplitudes [11477] = 8'd124;
   assign soundFileAmplitudes [11478] = 8'd132;
   assign soundFileAmplitudes [11479] = 8'd147;
   assign soundFileAmplitudes [11480] = 8'd145;
   assign soundFileAmplitudes [11481] = 8'd145;
   assign soundFileAmplitudes [11482] = 8'd142;
   assign soundFileAmplitudes [11483] = 8'd143;
   assign soundFileAmplitudes [11484] = 8'd144;
   assign soundFileAmplitudes [11485] = 8'd131;
   assign soundFileAmplitudes [11486] = 8'd125;
   assign soundFileAmplitudes [11487] = 8'd119;
   assign soundFileAmplitudes [11488] = 8'd104;
   assign soundFileAmplitudes [11489] = 8'd102;
   assign soundFileAmplitudes [11490] = 8'd113;
   assign soundFileAmplitudes [11491] = 8'd130;
   assign soundFileAmplitudes [11492] = 8'd132;
   assign soundFileAmplitudes [11493] = 8'd119;
   assign soundFileAmplitudes [11494] = 8'd108;
   assign soundFileAmplitudes [11495] = 8'd115;
   assign soundFileAmplitudes [11496] = 8'd122;
   assign soundFileAmplitudes [11497] = 8'd112;
   assign soundFileAmplitudes [11498] = 8'd109;
   assign soundFileAmplitudes [11499] = 8'd119;
   assign soundFileAmplitudes [11500] = 8'd130;
   assign soundFileAmplitudes [11501] = 8'd130;
   assign soundFileAmplitudes [11502] = 8'd104;
   assign soundFileAmplitudes [11503] = 8'd83;
   assign soundFileAmplitudes [11504] = 8'd96;
   assign soundFileAmplitudes [11505] = 8'd100;
   assign soundFileAmplitudes [11506] = 8'd123;
   assign soundFileAmplitudes [11507] = 8'd147;
   assign soundFileAmplitudes [11508] = 8'd140;
   assign soundFileAmplitudes [11509] = 8'd131;
   assign soundFileAmplitudes [11510] = 8'd133;
   assign soundFileAmplitudes [11511] = 8'd131;
   assign soundFileAmplitudes [11512] = 8'd153;
   assign soundFileAmplitudes [11513] = 8'd166;
   assign soundFileAmplitudes [11514] = 8'd160;
   assign soundFileAmplitudes [11515] = 8'd181;
   assign soundFileAmplitudes [11516] = 8'd172;
   assign soundFileAmplitudes [11517] = 8'd156;
   assign soundFileAmplitudes [11518] = 8'd143;
   assign soundFileAmplitudes [11519] = 8'd139;
   assign soundFileAmplitudes [11520] = 8'd126;
   assign soundFileAmplitudes [11521] = 8'd108;
   assign soundFileAmplitudes [11522] = 8'd107;
   assign soundFileAmplitudes [11523] = 8'd109;
   assign soundFileAmplitudes [11524] = 8'd111;
   assign soundFileAmplitudes [11525] = 8'd105;
   assign soundFileAmplitudes [11526] = 8'd96;
   assign soundFileAmplitudes [11527] = 8'd97;
   assign soundFileAmplitudes [11528] = 8'd116;
   assign soundFileAmplitudes [11529] = 8'd130;
   assign soundFileAmplitudes [11530] = 8'd128;
   assign soundFileAmplitudes [11531] = 8'd129;
   assign soundFileAmplitudes [11532] = 8'd125;
   assign soundFileAmplitudes [11533] = 8'd116;
   assign soundFileAmplitudes [11534] = 8'd109;
   assign soundFileAmplitudes [11535] = 8'd92;
   assign soundFileAmplitudes [11536] = 8'd96;
   assign soundFileAmplitudes [11537] = 8'd107;
   assign soundFileAmplitudes [11538] = 8'd113;
   assign soundFileAmplitudes [11539] = 8'd115;
   assign soundFileAmplitudes [11540] = 8'd110;
   assign soundFileAmplitudes [11541] = 8'd109;
   assign soundFileAmplitudes [11542] = 8'd114;
   assign soundFileAmplitudes [11543] = 8'd132;
   assign soundFileAmplitudes [11544] = 8'd149;
   assign soundFileAmplitudes [11545] = 8'd160;
   assign soundFileAmplitudes [11546] = 8'd151;
   assign soundFileAmplitudes [11547] = 8'd151;
   assign soundFileAmplitudes [11548] = 8'd157;
   assign soundFileAmplitudes [11549] = 8'd150;
   assign soundFileAmplitudes [11550] = 8'd156;
   assign soundFileAmplitudes [11551] = 8'd172;
   assign soundFileAmplitudes [11552] = 8'd165;
   assign soundFileAmplitudes [11553] = 8'd155;
   assign soundFileAmplitudes [11554] = 8'd151;
   assign soundFileAmplitudes [11555] = 8'd146;
   assign soundFileAmplitudes [11556] = 8'd134;
   assign soundFileAmplitudes [11557] = 8'd111;
   assign soundFileAmplitudes [11558] = 8'd107;
   assign soundFileAmplitudes [11559] = 8'd105;
   assign soundFileAmplitudes [11560] = 8'd114;
   assign soundFileAmplitudes [11561] = 8'd107;
   assign soundFileAmplitudes [11562] = 8'd97;
   assign soundFileAmplitudes [11563] = 8'd102;
   assign soundFileAmplitudes [11564] = 8'd109;
   assign soundFileAmplitudes [11565] = 8'd124;
   assign soundFileAmplitudes [11566] = 8'd111;
   assign soundFileAmplitudes [11567] = 8'd79;
   assign soundFileAmplitudes [11568] = 8'd79;
   assign soundFileAmplitudes [11569] = 8'd85;
   assign soundFileAmplitudes [11570] = 8'd94;
   assign soundFileAmplitudes [11571] = 8'd109;
   assign soundFileAmplitudes [11572] = 8'd110;
   assign soundFileAmplitudes [11573] = 8'd121;
   assign soundFileAmplitudes [11574] = 8'd132;
   assign soundFileAmplitudes [11575] = 8'd137;
   assign soundFileAmplitudes [11576] = 8'd157;
   assign soundFileAmplitudes [11577] = 8'd160;
   assign soundFileAmplitudes [11578] = 8'd149;
   assign soundFileAmplitudes [11579] = 8'd147;
   assign soundFileAmplitudes [11580] = 8'd149;
   assign soundFileAmplitudes [11581] = 8'd156;
   assign soundFileAmplitudes [11582] = 8'd153;
   assign soundFileAmplitudes [11583] = 8'd149;
   assign soundFileAmplitudes [11584] = 8'd146;
   assign soundFileAmplitudes [11585] = 8'd140;
   assign soundFileAmplitudes [11586] = 8'd133;
   assign soundFileAmplitudes [11587] = 8'd143;
   assign soundFileAmplitudes [11588] = 8'd148;
   assign soundFileAmplitudes [11589] = 8'd141;
   assign soundFileAmplitudes [11590] = 8'd133;
   assign soundFileAmplitudes [11591] = 8'd133;
   assign soundFileAmplitudes [11592] = 8'd133;
   assign soundFileAmplitudes [11593] = 8'd114;
   assign soundFileAmplitudes [11594] = 8'd107;
   assign soundFileAmplitudes [11595] = 8'd94;
   assign soundFileAmplitudes [11596] = 8'd102;
   assign soundFileAmplitudes [11597] = 8'd114;
   assign soundFileAmplitudes [11598] = 8'd100;
   assign soundFileAmplitudes [11599] = 8'd78;
   assign soundFileAmplitudes [11600] = 8'd64;
   assign soundFileAmplitudes [11601] = 8'd64;
   assign soundFileAmplitudes [11602] = 8'd75;
   assign soundFileAmplitudes [11603] = 8'd98;
   assign soundFileAmplitudes [11604] = 8'd104;
   assign soundFileAmplitudes [11605] = 8'd110;
   assign soundFileAmplitudes [11606] = 8'd119;
   assign soundFileAmplitudes [11607] = 8'd124;
   assign soundFileAmplitudes [11608] = 8'd131;
   assign soundFileAmplitudes [11609] = 8'd154;
   assign soundFileAmplitudes [11610] = 8'd176;
   assign soundFileAmplitudes [11611] = 8'd175;
   assign soundFileAmplitudes [11612] = 8'd166;
   assign soundFileAmplitudes [11613] = 8'd156;
   assign soundFileAmplitudes [11614] = 8'd150;
   assign soundFileAmplitudes [11615] = 8'd151;
   assign soundFileAmplitudes [11616] = 8'd149;
   assign soundFileAmplitudes [11617] = 8'd145;
   assign soundFileAmplitudes [11618] = 8'd147;
   assign soundFileAmplitudes [11619] = 8'd137;
   assign soundFileAmplitudes [11620] = 8'd126;
   assign soundFileAmplitudes [11621] = 8'd125;
   assign soundFileAmplitudes [11622] = 8'd118;
   assign soundFileAmplitudes [11623] = 8'd120;
   assign soundFileAmplitudes [11624] = 8'd127;
   assign soundFileAmplitudes [11625] = 8'd124;
   assign soundFileAmplitudes [11626] = 8'd124;
   assign soundFileAmplitudes [11627] = 8'd132;
   assign soundFileAmplitudes [11628] = 8'd132;
   assign soundFileAmplitudes [11629] = 8'd127;
   assign soundFileAmplitudes [11630] = 8'd126;
   assign soundFileAmplitudes [11631] = 8'd104;
   assign soundFileAmplitudes [11632] = 8'd80;
   assign soundFileAmplitudes [11633] = 8'd80;
   assign soundFileAmplitudes [11634] = 8'd86;
   assign soundFileAmplitudes [11635] = 8'd98;
   assign soundFileAmplitudes [11636] = 8'd99;
   assign soundFileAmplitudes [11637] = 8'd99;
   assign soundFileAmplitudes [11638] = 8'd100;
   assign soundFileAmplitudes [11639] = 8'd103;
   assign soundFileAmplitudes [11640] = 8'd104;
   assign soundFileAmplitudes [11641] = 8'd117;
   assign soundFileAmplitudes [11642] = 8'd145;
   assign soundFileAmplitudes [11643] = 8'd159;
   assign soundFileAmplitudes [11644] = 8'd160;
   assign soundFileAmplitudes [11645] = 8'd151;
   assign soundFileAmplitudes [11646] = 8'd149;
   assign soundFileAmplitudes [11647] = 8'd151;
   assign soundFileAmplitudes [11648] = 8'd161;
   assign soundFileAmplitudes [11649] = 8'd161;
   assign soundFileAmplitudes [11650] = 8'd151;
   assign soundFileAmplitudes [11651] = 8'd147;
   assign soundFileAmplitudes [11652] = 8'd142;
   assign soundFileAmplitudes [11653] = 8'd132;
   assign soundFileAmplitudes [11654] = 8'd118;
   assign soundFileAmplitudes [11655] = 8'd111;
   assign soundFileAmplitudes [11656] = 8'd116;
   assign soundFileAmplitudes [11657] = 8'd119;
   assign soundFileAmplitudes [11658] = 8'd123;
   assign soundFileAmplitudes [11659] = 8'd128;
   assign soundFileAmplitudes [11660] = 8'd153;
   assign soundFileAmplitudes [11661] = 8'd156;
   assign soundFileAmplitudes [11662] = 8'd149;
   assign soundFileAmplitudes [11663] = 8'd120;
   assign soundFileAmplitudes [11664] = 8'd83;
   assign soundFileAmplitudes [11665] = 8'd89;
   assign soundFileAmplitudes [11666] = 8'd97;
   assign soundFileAmplitudes [11667] = 8'd105;
   assign soundFileAmplitudes [11668] = 8'd102;
   assign soundFileAmplitudes [11669] = 8'd98;
   assign soundFileAmplitudes [11670] = 8'd94;
   assign soundFileAmplitudes [11671] = 8'd101;
   assign soundFileAmplitudes [11672] = 8'd108;
   assign soundFileAmplitudes [11673] = 8'd122;
   assign soundFileAmplitudes [11674] = 8'd135;
   assign soundFileAmplitudes [11675] = 8'd147;
   assign soundFileAmplitudes [11676] = 8'd144;
   assign soundFileAmplitudes [11677] = 8'd140;
   assign soundFileAmplitudes [11678] = 8'd134;
   assign soundFileAmplitudes [11679] = 8'd137;
   assign soundFileAmplitudes [11680] = 8'd156;
   assign soundFileAmplitudes [11681] = 8'd158;
   assign soundFileAmplitudes [11682] = 8'd152;
   assign soundFileAmplitudes [11683] = 8'd152;
   assign soundFileAmplitudes [11684] = 8'd155;
   assign soundFileAmplitudes [11685] = 8'd149;
   assign soundFileAmplitudes [11686] = 8'd144;
   assign soundFileAmplitudes [11687] = 8'd120;
   assign soundFileAmplitudes [11688] = 8'd111;
   assign soundFileAmplitudes [11689] = 8'd133;
   assign soundFileAmplitudes [11690] = 8'd146;
   assign soundFileAmplitudes [11691] = 8'd123;
   assign soundFileAmplitudes [11692] = 8'd115;
   assign soundFileAmplitudes [11693] = 8'd111;
   assign soundFileAmplitudes [11694] = 8'd111;
   assign soundFileAmplitudes [11695] = 8'd125;
   assign soundFileAmplitudes [11696] = 8'd110;
   assign soundFileAmplitudes [11697] = 8'd94;
   assign soundFileAmplitudes [11698] = 8'd87;
   assign soundFileAmplitudes [11699] = 8'd92;
   assign soundFileAmplitudes [11700] = 8'd104;
   assign soundFileAmplitudes [11701] = 8'd105;
   assign soundFileAmplitudes [11702] = 8'd90;
   assign soundFileAmplitudes [11703] = 8'd92;
   assign soundFileAmplitudes [11704] = 8'd95;
   assign soundFileAmplitudes [11705] = 8'd107;
   assign soundFileAmplitudes [11706] = 8'd122;
   assign soundFileAmplitudes [11707] = 8'd137;
   assign soundFileAmplitudes [11708] = 8'd156;
   assign soundFileAmplitudes [11709] = 8'd154;
   assign soundFileAmplitudes [11710] = 8'd154;
   assign soundFileAmplitudes [11711] = 8'd149;
   assign soundFileAmplitudes [11712] = 8'd154;
   assign soundFileAmplitudes [11713] = 8'd151;
   assign soundFileAmplitudes [11714] = 8'd138;
   assign soundFileAmplitudes [11715] = 8'd132;
   assign soundFileAmplitudes [11716] = 8'd139;
   assign soundFileAmplitudes [11717] = 8'd153;
   assign soundFileAmplitudes [11718] = 8'd150;
   assign soundFileAmplitudes [11719] = 8'd133;
   assign soundFileAmplitudes [11720] = 8'd123;
   assign soundFileAmplitudes [11721] = 8'd121;
   assign soundFileAmplitudes [11722] = 8'd117;
   assign soundFileAmplitudes [11723] = 8'd115;
   assign soundFileAmplitudes [11724] = 8'd110;
   assign soundFileAmplitudes [11725] = 8'd140;
   assign soundFileAmplitudes [11726] = 8'd153;
   assign soundFileAmplitudes [11727] = 8'd147;
   assign soundFileAmplitudes [11728] = 8'd148;
   assign soundFileAmplitudes [11729] = 8'd123;
   assign soundFileAmplitudes [11730] = 8'd96;
   assign soundFileAmplitudes [11731] = 8'd82;
   assign soundFileAmplitudes [11732] = 8'd92;
   assign soundFileAmplitudes [11733] = 8'd112;
   assign soundFileAmplitudes [11734] = 8'd120;
   assign soundFileAmplitudes [11735] = 8'd122;
   assign soundFileAmplitudes [11736] = 8'd123;
   assign soundFileAmplitudes [11737] = 8'd114;
   assign soundFileAmplitudes [11738] = 8'd109;
   assign soundFileAmplitudes [11739] = 8'd109;
   assign soundFileAmplitudes [11740] = 8'd124;
   assign soundFileAmplitudes [11741] = 8'd147;
   assign soundFileAmplitudes [11742] = 8'd142;
   assign soundFileAmplitudes [11743] = 8'd128;
   assign soundFileAmplitudes [11744] = 8'd123;
   assign soundFileAmplitudes [11745] = 8'd132;
   assign soundFileAmplitudes [11746] = 8'd141;
   assign soundFileAmplitudes [11747] = 8'd144;
   assign soundFileAmplitudes [11748] = 8'd152;
   assign soundFileAmplitudes [11749] = 8'd146;
   assign soundFileAmplitudes [11750] = 8'd139;
   assign soundFileAmplitudes [11751] = 8'd121;
   assign soundFileAmplitudes [11752] = 8'd100;
   assign soundFileAmplitudes [11753] = 8'd79;
   assign soundFileAmplitudes [11754] = 8'd87;
   assign soundFileAmplitudes [11755] = 8'd106;
   assign soundFileAmplitudes [11756] = 8'd121;
   assign soundFileAmplitudes [11757] = 8'd124;
   assign soundFileAmplitudes [11758] = 8'd103;
   assign soundFileAmplitudes [11759] = 8'd122;
   assign soundFileAmplitudes [11760] = 8'd133;
   assign soundFileAmplitudes [11761] = 8'd137;
   assign soundFileAmplitudes [11762] = 8'd120;
   assign soundFileAmplitudes [11763] = 8'd100;
   assign soundFileAmplitudes [11764] = 8'd116;
   assign soundFileAmplitudes [11765] = 8'd142;
   assign soundFileAmplitudes [11766] = 8'd160;
   assign soundFileAmplitudes [11767] = 8'd150;
   assign soundFileAmplitudes [11768] = 8'd136;
   assign soundFileAmplitudes [11769] = 8'd132;
   assign soundFileAmplitudes [11770] = 8'd128;
   assign soundFileAmplitudes [11771] = 8'd124;
   assign soundFileAmplitudes [11772] = 8'd129;
   assign soundFileAmplitudes [11773] = 8'd139;
   assign soundFileAmplitudes [11774] = 8'd140;
   assign soundFileAmplitudes [11775] = 8'd131;
   assign soundFileAmplitudes [11776] = 8'd129;
   assign soundFileAmplitudes [11777] = 8'd113;
   assign soundFileAmplitudes [11778] = 8'd107;
   assign soundFileAmplitudes [11779] = 8'd107;
   assign soundFileAmplitudes [11780] = 8'd115;
   assign soundFileAmplitudes [11781] = 8'd117;
   assign soundFileAmplitudes [11782] = 8'd131;
   assign soundFileAmplitudes [11783] = 8'd147;
   assign soundFileAmplitudes [11784] = 8'd139;
   assign soundFileAmplitudes [11785] = 8'd140;
   assign soundFileAmplitudes [11786] = 8'd134;
   assign soundFileAmplitudes [11787] = 8'd129;
   assign soundFileAmplitudes [11788] = 8'd128;
   assign soundFileAmplitudes [11789] = 8'd123;
   assign soundFileAmplitudes [11790] = 8'd114;
   assign soundFileAmplitudes [11791] = 8'd124;
   assign soundFileAmplitudes [11792] = 8'd126;
   assign soundFileAmplitudes [11793] = 8'd128;
   assign soundFileAmplitudes [11794] = 8'd115;
   assign soundFileAmplitudes [11795] = 8'd92;
   assign soundFileAmplitudes [11796] = 8'd99;
   assign soundFileAmplitudes [11797] = 8'd104;
   assign soundFileAmplitudes [11798] = 8'd119;
   assign soundFileAmplitudes [11799] = 8'd131;
   assign soundFileAmplitudes [11800] = 8'd135;
   assign soundFileAmplitudes [11801] = 8'd141;
   assign soundFileAmplitudes [11802] = 8'd151;
   assign soundFileAmplitudes [11803] = 8'd152;
   assign soundFileAmplitudes [11804] = 8'd162;
   assign soundFileAmplitudes [11805] = 8'd177;
   assign soundFileAmplitudes [11806] = 8'd166;
   assign soundFileAmplitudes [11807] = 8'd150;
   assign soundFileAmplitudes [11808] = 8'd141;
   assign soundFileAmplitudes [11809] = 8'd124;
   assign soundFileAmplitudes [11810] = 8'd113;
   assign soundFileAmplitudes [11811] = 8'd110;
   assign soundFileAmplitudes [11812] = 8'd110;
   assign soundFileAmplitudes [11813] = 8'd106;
   assign soundFileAmplitudes [11814] = 8'd93;
   assign soundFileAmplitudes [11815] = 8'd93;
   assign soundFileAmplitudes [11816] = 8'd88;
   assign soundFileAmplitudes [11817] = 8'd96;
   assign soundFileAmplitudes [11818] = 8'd105;
   assign soundFileAmplitudes [11819] = 8'd110;
   assign soundFileAmplitudes [11820] = 8'd117;
   assign soundFileAmplitudes [11821] = 8'd129;
   assign soundFileAmplitudes [11822] = 8'd131;
   assign soundFileAmplitudes [11823] = 8'd120;
   assign soundFileAmplitudes [11824] = 8'd128;
   assign soundFileAmplitudes [11825] = 8'd129;
   assign soundFileAmplitudes [11826] = 8'd142;
   assign soundFileAmplitudes [11827] = 8'd129;
   assign soundFileAmplitudes [11828] = 8'd104;
   assign soundFileAmplitudes [11829] = 8'd96;
   assign soundFileAmplitudes [11830] = 8'd94;
   assign soundFileAmplitudes [11831] = 8'd110;
   assign soundFileAmplitudes [11832] = 8'd124;
   assign soundFileAmplitudes [11833] = 8'd147;
   assign soundFileAmplitudes [11834] = 8'd147;
   assign soundFileAmplitudes [11835] = 8'd149;
   assign soundFileAmplitudes [11836] = 8'd163;
   assign soundFileAmplitudes [11837] = 8'd173;
   assign soundFileAmplitudes [11838] = 8'd182;
   assign soundFileAmplitudes [11839] = 8'd175;
   assign soundFileAmplitudes [11840] = 8'd175;
   assign soundFileAmplitudes [11841] = 8'd178;
   assign soundFileAmplitudes [11842] = 8'd171;
   assign soundFileAmplitudes [11843] = 8'd157;
   assign soundFileAmplitudes [11844] = 8'd139;
   assign soundFileAmplitudes [11845] = 8'd119;
   assign soundFileAmplitudes [11846] = 8'd93;
   assign soundFileAmplitudes [11847] = 8'd80;
   assign soundFileAmplitudes [11848] = 8'd83;
   assign soundFileAmplitudes [11849] = 8'd75;
   assign soundFileAmplitudes [11850] = 8'd74;
   assign soundFileAmplitudes [11851] = 8'd74;
   assign soundFileAmplitudes [11852] = 8'd73;
   assign soundFileAmplitudes [11853] = 8'd86;
   assign soundFileAmplitudes [11854] = 8'd97;
   assign soundFileAmplitudes [11855] = 8'd96;
   assign soundFileAmplitudes [11856] = 8'd105;
   assign soundFileAmplitudes [11857] = 8'd128;
   assign soundFileAmplitudes [11858] = 8'd125;
   assign soundFileAmplitudes [11859] = 8'd125;
   assign soundFileAmplitudes [11860] = 8'd100;
   assign soundFileAmplitudes [11861] = 8'd78;
   assign soundFileAmplitudes [11862] = 8'd99;
   assign soundFileAmplitudes [11863] = 8'd120;
   assign soundFileAmplitudes [11864] = 8'd142;
   assign soundFileAmplitudes [11865] = 8'd151;
   assign soundFileAmplitudes [11866] = 8'd152;
   assign soundFileAmplitudes [11867] = 8'd145;
   assign soundFileAmplitudes [11868] = 8'd157;
   assign soundFileAmplitudes [11869] = 8'd172;
   assign soundFileAmplitudes [11870] = 8'd176;
   assign soundFileAmplitudes [11871] = 8'd184;
   assign soundFileAmplitudes [11872] = 8'd183;
   assign soundFileAmplitudes [11873] = 8'd177;
   assign soundFileAmplitudes [11874] = 8'd178;
   assign soundFileAmplitudes [11875] = 8'd174;
   assign soundFileAmplitudes [11876] = 8'd154;
   assign soundFileAmplitudes [11877] = 8'd149;
   assign soundFileAmplitudes [11878] = 8'd142;
   assign soundFileAmplitudes [11879] = 8'd126;
   assign soundFileAmplitudes [11880] = 8'd127;
   assign soundFileAmplitudes [11881] = 8'd123;
   assign soundFileAmplitudes [11882] = 8'd95;
   assign soundFileAmplitudes [11883] = 8'd71;
   assign soundFileAmplitudes [11884] = 8'd53;
   assign soundFileAmplitudes [11885] = 8'd54;
   assign soundFileAmplitudes [11886] = 8'd60;
   assign soundFileAmplitudes [11887] = 8'd57;
   assign soundFileAmplitudes [11888] = 8'd62;
   assign soundFileAmplitudes [11889] = 8'd90;
   assign soundFileAmplitudes [11890] = 8'd108;
   assign soundFileAmplitudes [11891] = 8'd115;
   assign soundFileAmplitudes [11892] = 8'd110;
   assign soundFileAmplitudes [11893] = 8'd93;
   assign soundFileAmplitudes [11894] = 8'd92;
   assign soundFileAmplitudes [11895] = 8'd84;
   assign soundFileAmplitudes [11896] = 8'd108;
   assign soundFileAmplitudes [11897] = 8'd142;
   assign soundFileAmplitudes [11898] = 8'd157;
   assign soundFileAmplitudes [11899] = 8'd163;
   assign soundFileAmplitudes [11900] = 8'd163;
   assign soundFileAmplitudes [11901] = 8'd158;
   assign soundFileAmplitudes [11902] = 8'd167;
   assign soundFileAmplitudes [11903] = 8'd178;
   assign soundFileAmplitudes [11904] = 8'd185;
   assign soundFileAmplitudes [11905] = 8'd186;
   assign soundFileAmplitudes [11906] = 8'd180;
   assign soundFileAmplitudes [11907] = 8'd185;
   assign soundFileAmplitudes [11908] = 8'd175;
   assign soundFileAmplitudes [11909] = 8'd172;
   assign soundFileAmplitudes [11910] = 8'd165;
   assign soundFileAmplitudes [11911] = 8'd154;
   assign soundFileAmplitudes [11912] = 8'd144;
   assign soundFileAmplitudes [11913] = 8'd146;
   assign soundFileAmplitudes [11914] = 8'd134;
   assign soundFileAmplitudes [11915] = 8'd108;
   assign soundFileAmplitudes [11916] = 8'd89;
   assign soundFileAmplitudes [11917] = 8'd72;
   assign soundFileAmplitudes [11918] = 8'd80;
   assign soundFileAmplitudes [11919] = 8'd79;
   assign soundFileAmplitudes [11920] = 8'd71;
   assign soundFileAmplitudes [11921] = 8'd65;
   assign soundFileAmplitudes [11922] = 8'd73;
   assign soundFileAmplitudes [11923] = 8'd77;
   assign soundFileAmplitudes [11924] = 8'd79;
   assign soundFileAmplitudes [11925] = 8'd73;
   assign soundFileAmplitudes [11926] = 8'd71;
   assign soundFileAmplitudes [11927] = 8'd77;
   assign soundFileAmplitudes [11928] = 8'd88;
   assign soundFileAmplitudes [11929] = 8'd116;
   assign soundFileAmplitudes [11930] = 8'd129;
   assign soundFileAmplitudes [11931] = 8'd128;
   assign soundFileAmplitudes [11932] = 8'd116;
   assign soundFileAmplitudes [11933] = 8'd122;
   assign soundFileAmplitudes [11934] = 8'd144;
   assign soundFileAmplitudes [11935] = 8'd172;
   assign soundFileAmplitudes [11936] = 8'd184;
   assign soundFileAmplitudes [11937] = 8'd173;
   assign soundFileAmplitudes [11938] = 8'd161;
   assign soundFileAmplitudes [11939] = 8'd157;
   assign soundFileAmplitudes [11940] = 8'd176;
   assign soundFileAmplitudes [11941] = 8'd184;
   assign soundFileAmplitudes [11942] = 8'd177;
   assign soundFileAmplitudes [11943] = 8'd168;
   assign soundFileAmplitudes [11944] = 8'd169;
   assign soundFileAmplitudes [11945] = 8'd171;
   assign soundFileAmplitudes [11946] = 8'd164;
   assign soundFileAmplitudes [11947] = 8'd153;
   assign soundFileAmplitudes [11948] = 8'd141;
   assign soundFileAmplitudes [11949] = 8'd130;
   assign soundFileAmplitudes [11950] = 8'd111;
   assign soundFileAmplitudes [11951] = 8'd107;
   assign soundFileAmplitudes [11952] = 8'd108;
   assign soundFileAmplitudes [11953] = 8'd90;
   assign soundFileAmplitudes [11954] = 8'd86;
   assign soundFileAmplitudes [11955] = 8'd94;
   assign soundFileAmplitudes [11956] = 8'd87;
   assign soundFileAmplitudes [11957] = 8'd79;
   assign soundFileAmplitudes [11958] = 8'd56;
   assign soundFileAmplitudes [11959] = 8'd45;
   assign soundFileAmplitudes [11960] = 8'd59;
   assign soundFileAmplitudes [11961] = 8'd77;
   assign soundFileAmplitudes [11962] = 8'd103;
   assign soundFileAmplitudes [11963] = 8'd115;
   assign soundFileAmplitudes [11964] = 8'd127;
   assign soundFileAmplitudes [11965] = 8'd124;
   assign soundFileAmplitudes [11966] = 8'd131;
   assign soundFileAmplitudes [11967] = 8'd142;
   assign soundFileAmplitudes [11968] = 8'd146;
   assign soundFileAmplitudes [11969] = 8'd157;
   assign soundFileAmplitudes [11970] = 8'd151;
   assign soundFileAmplitudes [11971] = 8'd149;
   assign soundFileAmplitudes [11972] = 8'd154;
   assign soundFileAmplitudes [11973] = 8'd158;
   assign soundFileAmplitudes [11974] = 8'd147;
   assign soundFileAmplitudes [11975] = 8'd145;
   assign soundFileAmplitudes [11976] = 8'd162;
   assign soundFileAmplitudes [11977] = 8'd166;
   assign soundFileAmplitudes [11978] = 8'd168;
   assign soundFileAmplitudes [11979] = 8'd179;
   assign soundFileAmplitudes [11980] = 8'd167;
   assign soundFileAmplitudes [11981] = 8'd147;
   assign soundFileAmplitudes [11982] = 8'd133;
   assign soundFileAmplitudes [11983] = 8'd129;
   assign soundFileAmplitudes [11984] = 8'd129;
   assign soundFileAmplitudes [11985] = 8'd130;
   assign soundFileAmplitudes [11986] = 8'd129;
   assign soundFileAmplitudes [11987] = 8'd124;
   assign soundFileAmplitudes [11988] = 8'd120;
   assign soundFileAmplitudes [11989] = 8'd103;
   assign soundFileAmplitudes [11990] = 8'd86;
   assign soundFileAmplitudes [11991] = 8'd66;
   assign soundFileAmplitudes [11992] = 8'd61;
   assign soundFileAmplitudes [11993] = 8'd55;
   assign soundFileAmplitudes [11994] = 8'd58;
   assign soundFileAmplitudes [11995] = 8'd79;
   assign soundFileAmplitudes [11996] = 8'd92;
   assign soundFileAmplitudes [11997] = 8'd103;
   assign soundFileAmplitudes [11998] = 8'd107;
   assign soundFileAmplitudes [11999] = 8'd113;
   assign soundFileAmplitudes [12000] = 8'd121;
   assign soundFileAmplitudes [12001] = 8'd139;
   assign soundFileAmplitudes [12002] = 8'd153;
   assign soundFileAmplitudes [12003] = 8'd147;
   assign soundFileAmplitudes [12004] = 8'd139;
   assign soundFileAmplitudes [12005] = 8'd138;
   assign soundFileAmplitudes [12006] = 8'd152;
   assign soundFileAmplitudes [12007] = 8'd147;
   assign soundFileAmplitudes [12008] = 8'd134;
   assign soundFileAmplitudes [12009] = 8'd133;
   assign soundFileAmplitudes [12010] = 8'd135;
   assign soundFileAmplitudes [12011] = 8'd155;
   assign soundFileAmplitudes [12012] = 8'd158;
   assign soundFileAmplitudes [12013] = 8'd149;
   assign soundFileAmplitudes [12014] = 8'd142;
   assign soundFileAmplitudes [12015] = 8'd134;
   assign soundFileAmplitudes [12016] = 8'd137;
   assign soundFileAmplitudes [12017] = 8'd146;
   assign soundFileAmplitudes [12018] = 8'd147;
   assign soundFileAmplitudes [12019] = 8'd144;
   assign soundFileAmplitudes [12020] = 8'd154;
   assign soundFileAmplitudes [12021] = 8'd149;
   assign soundFileAmplitudes [12022] = 8'd142;
   assign soundFileAmplitudes [12023] = 8'd140;
   assign soundFileAmplitudes [12024] = 8'd123;
   assign soundFileAmplitudes [12025] = 8'd103;
   assign soundFileAmplitudes [12026] = 8'd91;
   assign soundFileAmplitudes [12027] = 8'd89;
   assign soundFileAmplitudes [12028] = 8'd91;
   assign soundFileAmplitudes [12029] = 8'd96;
   assign soundFileAmplitudes [12030] = 8'd84;
   assign soundFileAmplitudes [12031] = 8'd78;
   assign soundFileAmplitudes [12032] = 8'd89;
   assign soundFileAmplitudes [12033] = 8'd100;
   assign soundFileAmplitudes [12034] = 8'd110;
   assign soundFileAmplitudes [12035] = 8'd104;
   assign soundFileAmplitudes [12036] = 8'd114;
   assign soundFileAmplitudes [12037] = 8'd127;
   assign soundFileAmplitudes [12038] = 8'd133;
   assign soundFileAmplitudes [12039] = 8'd141;
   assign soundFileAmplitudes [12040] = 8'd138;
   assign soundFileAmplitudes [12041] = 8'd136;
   assign soundFileAmplitudes [12042] = 8'd148;
   assign soundFileAmplitudes [12043] = 8'd144;
   assign soundFileAmplitudes [12044] = 8'd143;
   assign soundFileAmplitudes [12045] = 8'd143;
   assign soundFileAmplitudes [12046] = 8'd133;
   assign soundFileAmplitudes [12047] = 8'd137;
   assign soundFileAmplitudes [12048] = 8'd134;
   assign soundFileAmplitudes [12049] = 8'd129;
   assign soundFileAmplitudes [12050] = 8'd134;
   assign soundFileAmplitudes [12051] = 8'd137;
   assign soundFileAmplitudes [12052] = 8'd129;
   assign soundFileAmplitudes [12053] = 8'd138;
   assign soundFileAmplitudes [12054] = 8'd149;
   assign soundFileAmplitudes [12055] = 8'd150;
   assign soundFileAmplitudes [12056] = 8'd148;
   assign soundFileAmplitudes [12057] = 8'd137;
   assign soundFileAmplitudes [12058] = 8'd131;
   assign soundFileAmplitudes [12059] = 8'd119;
   assign soundFileAmplitudes [12060] = 8'd106;
   assign soundFileAmplitudes [12061] = 8'd114;
   assign soundFileAmplitudes [12062] = 8'd126;
   assign soundFileAmplitudes [12063] = 8'd132;
   assign soundFileAmplitudes [12064] = 8'd128;
   assign soundFileAmplitudes [12065] = 8'd120;
   assign soundFileAmplitudes [12066] = 8'd104;
   assign soundFileAmplitudes [12067] = 8'd87;
   assign soundFileAmplitudes [12068] = 8'd94;
   assign soundFileAmplitudes [12069] = 8'd99;
   assign soundFileAmplitudes [12070] = 8'd104;
   assign soundFileAmplitudes [12071] = 8'd104;
   assign soundFileAmplitudes [12072] = 8'd111;
   assign soundFileAmplitudes [12073] = 8'd113;
   assign soundFileAmplitudes [12074] = 8'd115;
   assign soundFileAmplitudes [12075] = 8'd120;
   assign soundFileAmplitudes [12076] = 8'd120;
   assign soundFileAmplitudes [12077] = 8'd124;
   assign soundFileAmplitudes [12078] = 8'd137;
   assign soundFileAmplitudes [12079] = 8'd149;
   assign soundFileAmplitudes [12080] = 8'd142;
   assign soundFileAmplitudes [12081] = 8'd145;
   assign soundFileAmplitudes [12082] = 8'd137;
   assign soundFileAmplitudes [12083] = 8'd129;
   assign soundFileAmplitudes [12084] = 8'd126;
   assign soundFileAmplitudes [12085] = 8'd133;
   assign soundFileAmplitudes [12086] = 8'd144;
   assign soundFileAmplitudes [12087] = 8'd147;
   assign soundFileAmplitudes [12088] = 8'd150;
   assign soundFileAmplitudes [12089] = 8'd143;
   assign soundFileAmplitudes [12090] = 8'd145;
   assign soundFileAmplitudes [12091] = 8'd144;
   assign soundFileAmplitudes [12092] = 8'd126;
   assign soundFileAmplitudes [12093] = 8'd123;
   assign soundFileAmplitudes [12094] = 8'd128;
   assign soundFileAmplitudes [12095] = 8'd126;
   assign soundFileAmplitudes [12096] = 8'd133;
   assign soundFileAmplitudes [12097] = 8'd131;
   assign soundFileAmplitudes [12098] = 8'd126;
   assign soundFileAmplitudes [12099] = 8'd123;
   assign soundFileAmplitudes [12100] = 8'd116;
   assign soundFileAmplitudes [12101] = 8'd110;
   assign soundFileAmplitudes [12102] = 8'd106;
   assign soundFileAmplitudes [12103] = 8'd108;
   assign soundFileAmplitudes [12104] = 8'd116;
   assign soundFileAmplitudes [12105] = 8'd105;
   assign soundFileAmplitudes [12106] = 8'd103;
   assign soundFileAmplitudes [12107] = 8'd106;
   assign soundFileAmplitudes [12108] = 8'd103;
   assign soundFileAmplitudes [12109] = 8'd122;
   assign soundFileAmplitudes [12110] = 8'd144;
   assign soundFileAmplitudes [12111] = 8'd146;
   assign soundFileAmplitudes [12112] = 8'd138;
   assign soundFileAmplitudes [12113] = 8'd126;
   assign soundFileAmplitudes [12114] = 8'd121;
   assign soundFileAmplitudes [12115] = 8'd122;
   assign soundFileAmplitudes [12116] = 8'd121;
   assign soundFileAmplitudes [12117] = 8'd142;
   assign soundFileAmplitudes [12118] = 8'd144;
   assign soundFileAmplitudes [12119] = 8'd137;
   assign soundFileAmplitudes [12120] = 8'd135;
   assign soundFileAmplitudes [12121] = 8'd122;
   assign soundFileAmplitudes [12122] = 8'd120;
   assign soundFileAmplitudes [12123] = 8'd129;
   assign soundFileAmplitudes [12124] = 8'd130;
   assign soundFileAmplitudes [12125] = 8'd131;
   assign soundFileAmplitudes [12126] = 8'd127;
   assign soundFileAmplitudes [12127] = 8'd126;
   assign soundFileAmplitudes [12128] = 8'd130;
   assign soundFileAmplitudes [12129] = 8'd130;
   assign soundFileAmplitudes [12130] = 8'd131;
   assign soundFileAmplitudes [12131] = 8'd127;
   assign soundFileAmplitudes [12132] = 8'd127;
   assign soundFileAmplitudes [12133] = 8'd124;
   assign soundFileAmplitudes [12134] = 8'd127;
   assign soundFileAmplitudes [12135] = 8'd126;
   assign soundFileAmplitudes [12136] = 8'd115;
   assign soundFileAmplitudes [12137] = 8'd114;
   assign soundFileAmplitudes [12138] = 8'd112;
   assign soundFileAmplitudes [12139] = 8'd111;
   assign soundFileAmplitudes [12140] = 8'd125;
   assign soundFileAmplitudes [12141] = 8'd118;
   assign soundFileAmplitudes [12142] = 8'd118;
   assign soundFileAmplitudes [12143] = 8'd116;
   assign soundFileAmplitudes [12144] = 8'd110;
   assign soundFileAmplitudes [12145] = 8'd124;
   assign soundFileAmplitudes [12146] = 8'd136;
   assign soundFileAmplitudes [12147] = 8'd143;
   assign soundFileAmplitudes [12148] = 8'd133;
   assign soundFileAmplitudes [12149] = 8'd122;
   assign soundFileAmplitudes [12150] = 8'd118;
   assign soundFileAmplitudes [12151] = 8'd126;
   assign soundFileAmplitudes [12152] = 8'd130;
   assign soundFileAmplitudes [12153] = 8'd139;
   assign soundFileAmplitudes [12154] = 8'd127;
   assign soundFileAmplitudes [12155] = 8'd113;
   assign soundFileAmplitudes [12156] = 8'd115;
   assign soundFileAmplitudes [12157] = 8'd109;
   assign soundFileAmplitudes [12158] = 8'd116;
   assign soundFileAmplitudes [12159] = 8'd111;
   assign soundFileAmplitudes [12160] = 8'd107;
   assign soundFileAmplitudes [12161] = 8'd122;
   assign soundFileAmplitudes [12162] = 8'd133;
   assign soundFileAmplitudes [12163] = 8'd138;
   assign soundFileAmplitudes [12164] = 8'd143;
   assign soundFileAmplitudes [12165] = 8'd138;
   assign soundFileAmplitudes [12166] = 8'd130;
   assign soundFileAmplitudes [12167] = 8'd130;
   assign soundFileAmplitudes [12168] = 8'd137;
   assign soundFileAmplitudes [12169] = 8'd143;
   assign soundFileAmplitudes [12170] = 8'd144;
   assign soundFileAmplitudes [12171] = 8'd149;
   assign soundFileAmplitudes [12172] = 8'd142;
   assign soundFileAmplitudes [12173] = 8'd136;
   assign soundFileAmplitudes [12174] = 8'd124;
   assign soundFileAmplitudes [12175] = 8'd117;
   assign soundFileAmplitudes [12176] = 8'd121;
   assign soundFileAmplitudes [12177] = 8'd132;
   assign soundFileAmplitudes [12178] = 8'd126;
   assign soundFileAmplitudes [12179] = 8'd111;
   assign soundFileAmplitudes [12180] = 8'd112;
   assign soundFileAmplitudes [12181] = 8'd108;
   assign soundFileAmplitudes [12182] = 8'd114;
   assign soundFileAmplitudes [12183] = 8'd127;
   assign soundFileAmplitudes [12184] = 8'd127;
   assign soundFileAmplitudes [12185] = 8'd120;
   assign soundFileAmplitudes [12186] = 8'd116;
   assign soundFileAmplitudes [12187] = 8'd124;
   assign soundFileAmplitudes [12188] = 8'd136;
   assign soundFileAmplitudes [12189] = 8'd139;
   assign soundFileAmplitudes [12190] = 8'd136;
   assign soundFileAmplitudes [12191] = 8'd128;
   assign soundFileAmplitudes [12192] = 8'd121;
   assign soundFileAmplitudes [12193] = 8'd110;
   assign soundFileAmplitudes [12194] = 8'd99;
   assign soundFileAmplitudes [12195] = 8'd109;
   assign soundFileAmplitudes [12196] = 8'd121;
   assign soundFileAmplitudes [12197] = 8'd120;
   assign soundFileAmplitudes [12198] = 8'd125;
   assign soundFileAmplitudes [12199] = 8'd138;
   assign soundFileAmplitudes [12200] = 8'd145;
   assign soundFileAmplitudes [12201] = 8'd127;
   assign soundFileAmplitudes [12202] = 8'd118;
   assign soundFileAmplitudes [12203] = 8'd121;
   assign soundFileAmplitudes [12204] = 8'd127;
   assign soundFileAmplitudes [12205] = 8'd137;
   assign soundFileAmplitudes [12206] = 8'd139;
   assign soundFileAmplitudes [12207] = 8'd139;
   assign soundFileAmplitudes [12208] = 8'd140;
   assign soundFileAmplitudes [12209] = 8'd129;
   assign soundFileAmplitudes [12210] = 8'd114;
   assign soundFileAmplitudes [12211] = 8'd110;
   assign soundFileAmplitudes [12212] = 8'd112;
   assign soundFileAmplitudes [12213] = 8'd125;
   assign soundFileAmplitudes [12214] = 8'd122;
   assign soundFileAmplitudes [12215] = 8'd111;
   assign soundFileAmplitudes [12216] = 8'd104;
   assign soundFileAmplitudes [12217] = 8'd106;
   assign soundFileAmplitudes [12218] = 8'd116;
   assign soundFileAmplitudes [12219] = 8'd130;
   assign soundFileAmplitudes [12220] = 8'd135;
   assign soundFileAmplitudes [12221] = 8'd133;
   assign soundFileAmplitudes [12222] = 8'd128;
   assign soundFileAmplitudes [12223] = 8'd133;
   assign soundFileAmplitudes [12224] = 8'd152;
   assign soundFileAmplitudes [12225] = 8'd165;
   assign soundFileAmplitudes [12226] = 8'd167;
   assign soundFileAmplitudes [12227] = 8'd149;
   assign soundFileAmplitudes [12228] = 8'd133;
   assign soundFileAmplitudes [12229] = 8'd125;
   assign soundFileAmplitudes [12230] = 8'd114;
   assign soundFileAmplitudes [12231] = 8'd114;
   assign soundFileAmplitudes [12232] = 8'd114;
   assign soundFileAmplitudes [12233] = 8'd116;
   assign soundFileAmplitudes [12234] = 8'd114;
   assign soundFileAmplitudes [12235] = 8'd110;
   assign soundFileAmplitudes [12236] = 8'd118;
   assign soundFileAmplitudes [12237] = 8'd117;
   assign soundFileAmplitudes [12238] = 8'd122;
   assign soundFileAmplitudes [12239] = 8'd129;
   assign soundFileAmplitudes [12240] = 8'd134;
   assign soundFileAmplitudes [12241] = 8'd144;
   assign soundFileAmplitudes [12242] = 8'd147;
   assign soundFileAmplitudes [12243] = 8'd146;
   assign soundFileAmplitudes [12244] = 8'd140;
   assign soundFileAmplitudes [12245] = 8'd132;
   assign soundFileAmplitudes [12246] = 8'd127;
   assign soundFileAmplitudes [12247] = 8'd120;
   assign soundFileAmplitudes [12248] = 8'd117;
   assign soundFileAmplitudes [12249] = 8'd113;
   assign soundFileAmplitudes [12250] = 8'd102;
   assign soundFileAmplitudes [12251] = 8'd84;
   assign soundFileAmplitudes [12252] = 8'd78;
   assign soundFileAmplitudes [12253] = 8'd80;
   assign soundFileAmplitudes [12254] = 8'd98;
   assign soundFileAmplitudes [12255] = 8'd113;
   assign soundFileAmplitudes [12256] = 8'd116;
   assign soundFileAmplitudes [12257] = 8'd127;
   assign soundFileAmplitudes [12258] = 8'd130;
   assign soundFileAmplitudes [12259] = 8'd145;
   assign soundFileAmplitudes [12260] = 8'd157;
   assign soundFileAmplitudes [12261] = 8'd167;
   assign soundFileAmplitudes [12262] = 8'd171;
   assign soundFileAmplitudes [12263] = 8'd156;
   assign soundFileAmplitudes [12264] = 8'd146;
   assign soundFileAmplitudes [12265] = 8'd133;
   assign soundFileAmplitudes [12266] = 8'd122;
   assign soundFileAmplitudes [12267] = 8'd122;
   assign soundFileAmplitudes [12268] = 8'd129;
   assign soundFileAmplitudes [12269] = 8'd119;
   assign soundFileAmplitudes [12270] = 8'd107;
   assign soundFileAmplitudes [12271] = 8'd111;
   assign soundFileAmplitudes [12272] = 8'd116;
   assign soundFileAmplitudes [12273] = 8'd127;
   assign soundFileAmplitudes [12274] = 8'd132;
   assign soundFileAmplitudes [12275] = 8'd135;
   assign soundFileAmplitudes [12276] = 8'd128;
   assign soundFileAmplitudes [12277] = 8'd129;
   assign soundFileAmplitudes [12278] = 8'd144;
   assign soundFileAmplitudes [12279] = 8'd148;
   assign soundFileAmplitudes [12280] = 8'd142;
   assign soundFileAmplitudes [12281] = 8'd139;
   assign soundFileAmplitudes [12282] = 8'd136;
   assign soundFileAmplitudes [12283] = 8'd124;
   assign soundFileAmplitudes [12284] = 8'd113;
   assign soundFileAmplitudes [12285] = 8'd94;
   assign soundFileAmplitudes [12286] = 8'd84;
   assign soundFileAmplitudes [12287] = 8'd82;
   assign soundFileAmplitudes [12288] = 8'd76;
   assign soundFileAmplitudes [12289] = 8'd72;
   assign soundFileAmplitudes [12290] = 8'd80;
   assign soundFileAmplitudes [12291] = 8'd92;
   assign soundFileAmplitudes [12292] = 8'd111;
   assign soundFileAmplitudes [12293] = 8'd125;
   assign soundFileAmplitudes [12294] = 8'd135;
   assign soundFileAmplitudes [12295] = 8'd141;
   assign soundFileAmplitudes [12296] = 8'd164;
   assign soundFileAmplitudes [12297] = 8'd176;
   assign soundFileAmplitudes [12298] = 8'd172;
   assign soundFileAmplitudes [12299] = 8'd169;
   assign soundFileAmplitudes [12300] = 8'd153;
   assign soundFileAmplitudes [12301] = 8'd153;
   assign soundFileAmplitudes [12302] = 8'd138;
   assign soundFileAmplitudes [12303] = 8'd140;
   assign soundFileAmplitudes [12304] = 8'd149;
   assign soundFileAmplitudes [12305] = 8'd139;
   assign soundFileAmplitudes [12306] = 8'd131;
   assign soundFileAmplitudes [12307] = 8'd120;
   assign soundFileAmplitudes [12308] = 8'd109;
   assign soundFileAmplitudes [12309] = 8'd107;
   assign soundFileAmplitudes [12310] = 8'd118;
   assign soundFileAmplitudes [12311] = 8'd129;
   assign soundFileAmplitudes [12312] = 8'd124;
   assign soundFileAmplitudes [12313] = 8'd113;
   assign soundFileAmplitudes [12314] = 8'd113;
   assign soundFileAmplitudes [12315] = 8'd122;
   assign soundFileAmplitudes [12316] = 8'd132;
   assign soundFileAmplitudes [12317] = 8'd130;
   assign soundFileAmplitudes [12318] = 8'd126;
   assign soundFileAmplitudes [12319] = 8'd129;
   assign soundFileAmplitudes [12320] = 8'd121;
   assign soundFileAmplitudes [12321] = 8'd102;
   assign soundFileAmplitudes [12322] = 8'd81;
   assign soundFileAmplitudes [12323] = 8'd78;
   assign soundFileAmplitudes [12324] = 8'd82;
   assign soundFileAmplitudes [12325] = 8'd88;
   assign soundFileAmplitudes [12326] = 8'd98;
   assign soundFileAmplitudes [12327] = 8'd106;
   assign soundFileAmplitudes [12328] = 8'd117;
   assign soundFileAmplitudes [12329] = 8'd117;
   assign soundFileAmplitudes [12330] = 8'd122;
   assign soundFileAmplitudes [12331] = 8'd139;
   assign soundFileAmplitudes [12332] = 8'd158;
   assign soundFileAmplitudes [12333] = 8'd158;
   assign soundFileAmplitudes [12334] = 8'd170;
   assign soundFileAmplitudes [12335] = 8'd169;
   assign soundFileAmplitudes [12336] = 8'd154;
   assign soundFileAmplitudes [12337] = 8'd155;
   assign soundFileAmplitudes [12338] = 8'd143;
   assign soundFileAmplitudes [12339] = 8'd139;
   assign soundFileAmplitudes [12340] = 8'd137;
   assign soundFileAmplitudes [12341] = 8'd146;
   assign soundFileAmplitudes [12342] = 8'd159;
   assign soundFileAmplitudes [12343] = 8'd153;
   assign soundFileAmplitudes [12344] = 8'd133;
   assign soundFileAmplitudes [12345] = 8'd111;
   assign soundFileAmplitudes [12346] = 8'd104;
   assign soundFileAmplitudes [12347] = 8'd115;
   assign soundFileAmplitudes [12348] = 8'd135;
   assign soundFileAmplitudes [12349] = 8'd147;
   assign soundFileAmplitudes [12350] = 8'd140;
   assign soundFileAmplitudes [12351] = 8'd117;
   assign soundFileAmplitudes [12352] = 8'd106;
   assign soundFileAmplitudes [12353] = 8'd119;
   assign soundFileAmplitudes [12354] = 8'd123;
   assign soundFileAmplitudes [12355] = 8'd122;
   assign soundFileAmplitudes [12356] = 8'd124;
   assign soundFileAmplitudes [12357] = 8'd108;
   assign soundFileAmplitudes [12358] = 8'd85;
   assign soundFileAmplitudes [12359] = 8'd66;
   assign soundFileAmplitudes [12360] = 8'd61;
   assign soundFileAmplitudes [12361] = 8'd72;
   assign soundFileAmplitudes [12362] = 8'd92;
   assign soundFileAmplitudes [12363] = 8'd113;
   assign soundFileAmplitudes [12364] = 8'd116;
   assign soundFileAmplitudes [12365] = 8'd110;
   assign soundFileAmplitudes [12366] = 8'd104;
   assign soundFileAmplitudes [12367] = 8'd111;
   assign soundFileAmplitudes [12368] = 8'd149;
   assign soundFileAmplitudes [12369] = 8'd164;
   assign soundFileAmplitudes [12370] = 8'd177;
   assign soundFileAmplitudes [12371] = 8'd177;
   assign soundFileAmplitudes [12372] = 8'd161;
   assign soundFileAmplitudes [12373] = 8'd164;
   assign soundFileAmplitudes [12374] = 8'd168;
   assign soundFileAmplitudes [12375] = 8'd168;
   assign soundFileAmplitudes [12376] = 8'd167;
   assign soundFileAmplitudes [12377] = 8'd156;
   assign soundFileAmplitudes [12378] = 8'd143;
   assign soundFileAmplitudes [12379] = 8'd142;
   assign soundFileAmplitudes [12380] = 8'd133;
   assign soundFileAmplitudes [12381] = 8'd128;
   assign soundFileAmplitudes [12382] = 8'd110;
   assign soundFileAmplitudes [12383] = 8'd98;
   assign soundFileAmplitudes [12384] = 8'd89;
   assign soundFileAmplitudes [12385] = 8'd87;
   assign soundFileAmplitudes [12386] = 8'd103;
   assign soundFileAmplitudes [12387] = 8'd113;
   assign soundFileAmplitudes [12388] = 8'd121;
   assign soundFileAmplitudes [12389] = 8'd121;
   assign soundFileAmplitudes [12390] = 8'd123;
   assign soundFileAmplitudes [12391] = 8'd124;
   assign soundFileAmplitudes [12392] = 8'd132;
   assign soundFileAmplitudes [12393] = 8'd140;
   assign soundFileAmplitudes [12394] = 8'd126;
   assign soundFileAmplitudes [12395] = 8'd101;
   assign soundFileAmplitudes [12396] = 8'd84;
   assign soundFileAmplitudes [12397] = 8'd82;
   assign soundFileAmplitudes [12398] = 8'd86;
   assign soundFileAmplitudes [12399] = 8'd104;
   assign soundFileAmplitudes [12400] = 8'd115;
   assign soundFileAmplitudes [12401] = 8'd115;
   assign soundFileAmplitudes [12402] = 8'd111;
   assign soundFileAmplitudes [12403] = 8'd108;
   assign soundFileAmplitudes [12404] = 8'd124;
   assign soundFileAmplitudes [12405] = 8'd127;
   assign soundFileAmplitudes [12406] = 8'd140;
   assign soundFileAmplitudes [12407] = 8'd152;
   assign soundFileAmplitudes [12408] = 8'd160;
   assign soundFileAmplitudes [12409] = 8'd171;
   assign soundFileAmplitudes [12410] = 8'd167;
   assign soundFileAmplitudes [12411] = 8'd160;
   assign soundFileAmplitudes [12412] = 8'd161;
   assign soundFileAmplitudes [12413] = 8'd163;
   assign soundFileAmplitudes [12414] = 8'd155;
   assign soundFileAmplitudes [12415] = 8'd142;
   assign soundFileAmplitudes [12416] = 8'd129;
   assign soundFileAmplitudes [12417] = 8'd120;
   assign soundFileAmplitudes [12418] = 8'd105;
   assign soundFileAmplitudes [12419] = 8'd99;
   assign soundFileAmplitudes [12420] = 8'd94;
   assign soundFileAmplitudes [12421] = 8'd102;
   assign soundFileAmplitudes [12422] = 8'd114;
   assign soundFileAmplitudes [12423] = 8'd119;
   assign soundFileAmplitudes [12424] = 8'd135;
   assign soundFileAmplitudes [12425] = 8'd133;
   assign soundFileAmplitudes [12426] = 8'd132;
   assign soundFileAmplitudes [12427] = 8'd123;
   assign soundFileAmplitudes [12428] = 8'd135;
   assign soundFileAmplitudes [12429] = 8'd145;
   assign soundFileAmplitudes [12430] = 8'd157;
   assign soundFileAmplitudes [12431] = 8'd145;
   assign soundFileAmplitudes [12432] = 8'd93;
   assign soundFileAmplitudes [12433] = 8'd91;
   assign soundFileAmplitudes [12434] = 8'd83;
   assign soundFileAmplitudes [12435] = 8'd85;
   assign soundFileAmplitudes [12436] = 8'd97;
   assign soundFileAmplitudes [12437] = 8'd94;
   assign soundFileAmplitudes [12438] = 8'd87;
   assign soundFileAmplitudes [12439] = 8'd110;
   assign soundFileAmplitudes [12440] = 8'd128;
   assign soundFileAmplitudes [12441] = 8'd128;
   assign soundFileAmplitudes [12442] = 8'd128;
   assign soundFileAmplitudes [12443] = 8'd116;
   assign soundFileAmplitudes [12444] = 8'd131;
   assign soundFileAmplitudes [12445] = 8'd149;
   assign soundFileAmplitudes [12446] = 8'd158;
   assign soundFileAmplitudes [12447] = 8'd164;
   assign soundFileAmplitudes [12448] = 8'd155;
   assign soundFileAmplitudes [12449] = 8'd150;
   assign soundFileAmplitudes [12450] = 8'd149;
   assign soundFileAmplitudes [12451] = 8'd152;
   assign soundFileAmplitudes [12452] = 8'd156;
   assign soundFileAmplitudes [12453] = 8'd148;
   assign soundFileAmplitudes [12454] = 8'd138;
   assign soundFileAmplitudes [12455] = 8'd125;
   assign soundFileAmplitudes [12456] = 8'd116;
   assign soundFileAmplitudes [12457] = 8'd111;
   assign soundFileAmplitudes [12458] = 8'd116;
   assign soundFileAmplitudes [12459] = 8'd111;
   assign soundFileAmplitudes [12460] = 8'd119;
   assign soundFileAmplitudes [12461] = 8'd129;
   assign soundFileAmplitudes [12462] = 8'd129;
   assign soundFileAmplitudes [12463] = 8'd130;
   assign soundFileAmplitudes [12464] = 8'd132;
   assign soundFileAmplitudes [12465] = 8'd140;
   assign soundFileAmplitudes [12466] = 8'd133;
   assign soundFileAmplitudes [12467] = 8'd118;
   assign soundFileAmplitudes [12468] = 8'd103;
   assign soundFileAmplitudes [12469] = 8'd90;
   assign soundFileAmplitudes [12470] = 8'd83;
   assign soundFileAmplitudes [12471] = 8'd89;
   assign soundFileAmplitudes [12472] = 8'd96;
   assign soundFileAmplitudes [12473] = 8'd108;
   assign soundFileAmplitudes [12474] = 8'd117;
   assign soundFileAmplitudes [12475] = 8'd123;
   assign soundFileAmplitudes [12476] = 8'd123;
   assign soundFileAmplitudes [12477] = 8'd127;
   assign soundFileAmplitudes [12478] = 8'd130;
   assign soundFileAmplitudes [12479] = 8'd124;
   assign soundFileAmplitudes [12480] = 8'd120;
   assign soundFileAmplitudes [12481] = 8'd129;
   assign soundFileAmplitudes [12482] = 8'd140;
   assign soundFileAmplitudes [12483] = 8'd151;
   assign soundFileAmplitudes [12484] = 8'd144;
   assign soundFileAmplitudes [12485] = 8'd136;
   assign soundFileAmplitudes [12486] = 8'd138;
   assign soundFileAmplitudes [12487] = 8'd130;
   assign soundFileAmplitudes [12488] = 8'd147;
   assign soundFileAmplitudes [12489] = 8'd144;
   assign soundFileAmplitudes [12490] = 8'd147;
   assign soundFileAmplitudes [12491] = 8'd137;
   assign soundFileAmplitudes [12492] = 8'd116;
   assign soundFileAmplitudes [12493] = 8'd118;
   assign soundFileAmplitudes [12494] = 8'd127;
   assign soundFileAmplitudes [12495] = 8'd132;
   assign soundFileAmplitudes [12496] = 8'd126;
   assign soundFileAmplitudes [12497] = 8'd132;
   assign soundFileAmplitudes [12498] = 8'd127;
   assign soundFileAmplitudes [12499] = 8'd119;
   assign soundFileAmplitudes [12500] = 8'd114;
   assign soundFileAmplitudes [12501] = 8'd129;
   assign soundFileAmplitudes [12502] = 8'd132;
   assign soundFileAmplitudes [12503] = 8'd130;
   assign soundFileAmplitudes [12504] = 8'd134;
   assign soundFileAmplitudes [12505] = 8'd120;
   assign soundFileAmplitudes [12506] = 8'd115;
   assign soundFileAmplitudes [12507] = 8'd111;
   assign soundFileAmplitudes [12508] = 8'd99;
   assign soundFileAmplitudes [12509] = 8'd98;
   assign soundFileAmplitudes [12510] = 8'd113;
   assign soundFileAmplitudes [12511] = 8'd117;
   assign soundFileAmplitudes [12512] = 8'd115;
   assign soundFileAmplitudes [12513] = 8'd131;
   assign soundFileAmplitudes [12514] = 8'd133;
   assign soundFileAmplitudes [12515] = 8'd118;
   assign soundFileAmplitudes [12516] = 8'd128;
   assign soundFileAmplitudes [12517] = 8'd121;
   assign soundFileAmplitudes [12518] = 8'd133;
   assign soundFileAmplitudes [12519] = 8'd144;
   assign soundFileAmplitudes [12520] = 8'd148;
   assign soundFileAmplitudes [12521] = 8'd150;
   assign soundFileAmplitudes [12522] = 8'd138;
   assign soundFileAmplitudes [12523] = 8'd127;
   assign soundFileAmplitudes [12524] = 8'd118;
   assign soundFileAmplitudes [12525] = 8'd128;
   assign soundFileAmplitudes [12526] = 8'd134;
   assign soundFileAmplitudes [12527] = 8'd148;
   assign soundFileAmplitudes [12528] = 8'd137;
   assign soundFileAmplitudes [12529] = 8'd129;
   assign soundFileAmplitudes [12530] = 8'd128;
   assign soundFileAmplitudes [12531] = 8'd126;
   assign soundFileAmplitudes [12532] = 8'd121;
   assign soundFileAmplitudes [12533] = 8'd115;
   assign soundFileAmplitudes [12534] = 8'd110;
   assign soundFileAmplitudes [12535] = 8'd104;
   assign soundFileAmplitudes [12536] = 8'd101;
   assign soundFileAmplitudes [12537] = 8'd115;
   assign soundFileAmplitudes [12538] = 8'd128;
   assign soundFileAmplitudes [12539] = 8'd130;
   assign soundFileAmplitudes [12540] = 8'd145;
   assign soundFileAmplitudes [12541] = 8'd136;
   assign soundFileAmplitudes [12542] = 8'd123;
   assign soundFileAmplitudes [12543] = 8'd116;
   assign soundFileAmplitudes [12544] = 8'd100;
   assign soundFileAmplitudes [12545] = 8'd94;
   assign soundFileAmplitudes [12546] = 8'd101;
   assign soundFileAmplitudes [12547] = 8'd118;
   assign soundFileAmplitudes [12548] = 8'd126;
   assign soundFileAmplitudes [12549] = 8'd112;
   assign soundFileAmplitudes [12550] = 8'd121;
   assign soundFileAmplitudes [12551] = 8'd125;
   assign soundFileAmplitudes [12552] = 8'd134;
   assign soundFileAmplitudes [12553] = 8'd138;
   assign soundFileAmplitudes [12554] = 8'd123;
   assign soundFileAmplitudes [12555] = 8'd131;
   assign soundFileAmplitudes [12556] = 8'd146;
   assign soundFileAmplitudes [12557] = 8'd146;
   assign soundFileAmplitudes [12558] = 8'd139;
   assign soundFileAmplitudes [12559] = 8'd133;
   assign soundFileAmplitudes [12560] = 8'd129;
   assign soundFileAmplitudes [12561] = 8'd131;
   assign soundFileAmplitudes [12562] = 8'd135;
   assign soundFileAmplitudes [12563] = 8'd153;
   assign soundFileAmplitudes [12564] = 8'd148;
   assign soundFileAmplitudes [12565] = 8'd135;
   assign soundFileAmplitudes [12566] = 8'd128;
   assign soundFileAmplitudes [12567] = 8'd121;
   assign soundFileAmplitudes [12568] = 8'd130;
   assign soundFileAmplitudes [12569] = 8'd135;
   assign soundFileAmplitudes [12570] = 8'd133;
   assign soundFileAmplitudes [12571] = 8'd128;
   assign soundFileAmplitudes [12572] = 8'd112;
   assign soundFileAmplitudes [12573] = 8'd101;
   assign soundFileAmplitudes [12574] = 8'd109;
   assign soundFileAmplitudes [12575] = 8'd116;
   assign soundFileAmplitudes [12576] = 8'd122;
   assign soundFileAmplitudes [12577] = 8'd128;
   assign soundFileAmplitudes [12578] = 8'd127;
   assign soundFileAmplitudes [12579] = 8'd123;
   assign soundFileAmplitudes [12580] = 8'd107;
   assign soundFileAmplitudes [12581] = 8'd107;
   assign soundFileAmplitudes [12582] = 8'd110;
   assign soundFileAmplitudes [12583] = 8'd113;
   assign soundFileAmplitudes [12584] = 8'd124;
   assign soundFileAmplitudes [12585] = 8'd130;
   assign soundFileAmplitudes [12586] = 8'd124;
   assign soundFileAmplitudes [12587] = 8'd113;
   assign soundFileAmplitudes [12588] = 8'd115;
   assign soundFileAmplitudes [12589] = 8'd126;
   assign soundFileAmplitudes [12590] = 8'd138;
   assign soundFileAmplitudes [12591] = 8'd120;
   assign soundFileAmplitudes [12592] = 8'd115;
   assign soundFileAmplitudes [12593] = 8'd135;
   assign soundFileAmplitudes [12594] = 8'd133;
   assign soundFileAmplitudes [12595] = 8'd132;
   assign soundFileAmplitudes [12596] = 8'd136;
   assign soundFileAmplitudes [12597] = 8'd134;
   assign soundFileAmplitudes [12598] = 8'd121;
   assign soundFileAmplitudes [12599] = 8'd131;
   assign soundFileAmplitudes [12600] = 8'd140;
   assign soundFileAmplitudes [12601] = 8'd138;
   assign soundFileAmplitudes [12602] = 8'd141;
   assign soundFileAmplitudes [12603] = 8'd137;
   assign soundFileAmplitudes [12604] = 8'd135;
   assign soundFileAmplitudes [12605] = 8'd130;
   assign soundFileAmplitudes [12606] = 8'd137;
   assign soundFileAmplitudes [12607] = 8'd130;
   assign soundFileAmplitudes [12608] = 8'd120;
   assign soundFileAmplitudes [12609] = 8'd124;
   assign soundFileAmplitudes [12610] = 8'd131;
   assign soundFileAmplitudes [12611] = 8'd105;
   assign soundFileAmplitudes [12612] = 8'd105;
   assign soundFileAmplitudes [12613] = 8'd112;
   assign soundFileAmplitudes [12614] = 8'd122;
   assign soundFileAmplitudes [12615] = 8'd140;
   assign soundFileAmplitudes [12616] = 8'd136;
   assign soundFileAmplitudes [12617] = 8'd121;
   assign soundFileAmplitudes [12618] = 8'd113;
   assign soundFileAmplitudes [12619] = 8'd112;
   assign soundFileAmplitudes [12620] = 8'd108;
   assign soundFileAmplitudes [12621] = 8'd124;
   assign soundFileAmplitudes [12622] = 8'd129;
   assign soundFileAmplitudes [12623] = 8'd126;
   assign soundFileAmplitudes [12624] = 8'd98;
   assign soundFileAmplitudes [12625] = 8'd123;
   assign soundFileAmplitudes [12626] = 8'd128;
   assign soundFileAmplitudes [12627] = 8'd135;
   assign soundFileAmplitudes [12628] = 8'd134;
   assign soundFileAmplitudes [12629] = 8'd119;
   assign soundFileAmplitudes [12630] = 8'd134;
   assign soundFileAmplitudes [12631] = 8'd124;
   assign soundFileAmplitudes [12632] = 8'd124;
   assign soundFileAmplitudes [12633] = 8'd131;
   assign soundFileAmplitudes [12634] = 8'd137;
   assign soundFileAmplitudes [12635] = 8'd125;
   assign soundFileAmplitudes [12636] = 8'd129;
   assign soundFileAmplitudes [12637] = 8'd134;
   assign soundFileAmplitudes [12638] = 8'd135;
   assign soundFileAmplitudes [12639] = 8'd134;
   assign soundFileAmplitudes [12640] = 8'd140;
   assign soundFileAmplitudes [12641] = 8'd138;
   assign soundFileAmplitudes [12642] = 8'd146;
   assign soundFileAmplitudes [12643] = 8'd140;
   assign soundFileAmplitudes [12644] = 8'd122;
   assign soundFileAmplitudes [12645] = 8'd116;
   assign soundFileAmplitudes [12646] = 8'd131;
   assign soundFileAmplitudes [12647] = 8'd131;
   assign soundFileAmplitudes [12648] = 8'd115;
   assign soundFileAmplitudes [12649] = 8'd109;
   assign soundFileAmplitudes [12650] = 8'd107;
   assign soundFileAmplitudes [12651] = 8'd121;
   assign soundFileAmplitudes [12652] = 8'd120;
   assign soundFileAmplitudes [12653] = 8'd125;
   assign soundFileAmplitudes [12654] = 8'd122;
   assign soundFileAmplitudes [12655] = 8'd118;
   assign soundFileAmplitudes [12656] = 8'd127;
   assign soundFileAmplitudes [12657] = 8'd130;
   assign soundFileAmplitudes [12658] = 8'd109;
   assign soundFileAmplitudes [12659] = 8'd122;
   assign soundFileAmplitudes [12660] = 8'd120;
   assign soundFileAmplitudes [12661] = 8'd129;
   assign soundFileAmplitudes [12662] = 8'd128;
   assign soundFileAmplitudes [12663] = 8'd124;
   assign soundFileAmplitudes [12664] = 8'd135;
   assign soundFileAmplitudes [12665] = 8'd129;
   assign soundFileAmplitudes [12666] = 8'd131;
   assign soundFileAmplitudes [12667] = 8'd109;
   assign soundFileAmplitudes [12668] = 8'd110;
   assign soundFileAmplitudes [12669] = 8'd107;
   assign soundFileAmplitudes [12670] = 8'd105;
   assign soundFileAmplitudes [12671] = 8'd111;
   assign soundFileAmplitudes [12672] = 8'd124;
   assign soundFileAmplitudes [12673] = 8'd116;
   assign soundFileAmplitudes [12674] = 8'd119;
   assign soundFileAmplitudes [12675] = 8'd135;
   assign soundFileAmplitudes [12676] = 8'd150;
   assign soundFileAmplitudes [12677] = 8'd156;
   assign soundFileAmplitudes [12678] = 8'd147;
   assign soundFileAmplitudes [12679] = 8'd147;
   assign soundFileAmplitudes [12680] = 8'd143;
   assign soundFileAmplitudes [12681] = 8'd138;
   assign soundFileAmplitudes [12682] = 8'd147;
   assign soundFileAmplitudes [12683] = 8'd141;
   assign soundFileAmplitudes [12684] = 8'd123;
   assign soundFileAmplitudes [12685] = 8'd113;
   assign soundFileAmplitudes [12686] = 8'd93;
   assign soundFileAmplitudes [12687] = 8'd94;
   assign soundFileAmplitudes [12688] = 8'd109;
   assign soundFileAmplitudes [12689] = 8'd126;
   assign soundFileAmplitudes [12690] = 8'd132;
   assign soundFileAmplitudes [12691] = 8'd135;
   assign soundFileAmplitudes [12692] = 8'd124;
   assign soundFileAmplitudes [12693] = 8'd123;
   assign soundFileAmplitudes [12694] = 8'd124;
   assign soundFileAmplitudes [12695] = 8'd127;
   assign soundFileAmplitudes [12696] = 8'd118;
   assign soundFileAmplitudes [12697] = 8'd105;
   assign soundFileAmplitudes [12698] = 8'd122;
   assign soundFileAmplitudes [12699] = 8'd125;
   assign soundFileAmplitudes [12700] = 8'd118;
   assign soundFileAmplitudes [12701] = 8'd130;
   assign soundFileAmplitudes [12702] = 8'd127;
   assign soundFileAmplitudes [12703] = 8'd114;
   assign soundFileAmplitudes [12704] = 8'd110;
   assign soundFileAmplitudes [12705] = 8'd96;
   assign soundFileAmplitudes [12706] = 8'd114;
   assign soundFileAmplitudes [12707] = 8'd117;
   assign soundFileAmplitudes [12708] = 8'd130;
   assign soundFileAmplitudes [12709] = 8'd135;
   assign soundFileAmplitudes [12710] = 8'd126;
   assign soundFileAmplitudes [12711] = 8'd133;
   assign soundFileAmplitudes [12712] = 8'd154;
   assign soundFileAmplitudes [12713] = 8'd169;
   assign soundFileAmplitudes [12714] = 8'd171;
   assign soundFileAmplitudes [12715] = 8'd162;
   assign soundFileAmplitudes [12716] = 8'd143;
   assign soundFileAmplitudes [12717] = 8'd137;
   assign soundFileAmplitudes [12718] = 8'd135;
   assign soundFileAmplitudes [12719] = 8'd143;
   assign soundFileAmplitudes [12720] = 8'd125;
   assign soundFileAmplitudes [12721] = 8'd120;
   assign soundFileAmplitudes [12722] = 8'd121;
   assign soundFileAmplitudes [12723] = 8'd115;
   assign soundFileAmplitudes [12724] = 8'd106;
   assign soundFileAmplitudes [12725] = 8'd89;
   assign soundFileAmplitudes [12726] = 8'd98;
   assign soundFileAmplitudes [12727] = 8'd105;
   assign soundFileAmplitudes [12728] = 8'd115;
   assign soundFileAmplitudes [12729] = 8'd123;
   assign soundFileAmplitudes [12730] = 8'd114;
   assign soundFileAmplitudes [12731] = 8'd120;
   assign soundFileAmplitudes [12732] = 8'd108;
   assign soundFileAmplitudes [12733] = 8'd109;
   assign soundFileAmplitudes [12734] = 8'd121;
   assign soundFileAmplitudes [12735] = 8'd121;
   assign soundFileAmplitudes [12736] = 8'd119;
   assign soundFileAmplitudes [12737] = 8'd128;
   assign soundFileAmplitudes [12738] = 8'd125;
   assign soundFileAmplitudes [12739] = 8'd126;
   assign soundFileAmplitudes [12740] = 8'd149;
   assign soundFileAmplitudes [12741] = 8'd154;
   assign soundFileAmplitudes [12742] = 8'd154;
   assign soundFileAmplitudes [12743] = 8'd119;
   assign soundFileAmplitudes [12744] = 8'd127;
   assign soundFileAmplitudes [12745] = 8'd135;
   assign soundFileAmplitudes [12746] = 8'd132;
   assign soundFileAmplitudes [12747] = 8'd138;
   assign soundFileAmplitudes [12748] = 8'd125;
   assign soundFileAmplitudes [12749] = 8'd131;
   assign soundFileAmplitudes [12750] = 8'd142;
   assign soundFileAmplitudes [12751] = 8'd152;
   assign soundFileAmplitudes [12752] = 8'd149;
   assign soundFileAmplitudes [12753] = 8'd135;
   assign soundFileAmplitudes [12754] = 8'd131;
   assign soundFileAmplitudes [12755] = 8'd140;
   assign soundFileAmplitudes [12756] = 8'd125;
   assign soundFileAmplitudes [12757] = 8'd104;
   assign soundFileAmplitudes [12758] = 8'd105;
   assign soundFileAmplitudes [12759] = 8'd111;
   assign soundFileAmplitudes [12760] = 8'd112;
   assign soundFileAmplitudes [12761] = 8'd99;
   assign soundFileAmplitudes [12762] = 8'd89;
   assign soundFileAmplitudes [12763] = 8'd91;
   assign soundFileAmplitudes [12764] = 8'd107;
   assign soundFileAmplitudes [12765] = 8'd128;
   assign soundFileAmplitudes [12766] = 8'd130;
   assign soundFileAmplitudes [12767] = 8'd127;
   assign soundFileAmplitudes [12768] = 8'd106;
   assign soundFileAmplitudes [12769] = 8'd108;
   assign soundFileAmplitudes [12770] = 8'd131;
   assign soundFileAmplitudes [12771] = 8'd135;
   assign soundFileAmplitudes [12772] = 8'd138;
   assign soundFileAmplitudes [12773] = 8'd139;
   assign soundFileAmplitudes [12774] = 8'd139;
   assign soundFileAmplitudes [12775] = 8'd138;
   assign soundFileAmplitudes [12776] = 8'd140;
   assign soundFileAmplitudes [12777] = 8'd137;
   assign soundFileAmplitudes [12778] = 8'd126;
   assign soundFileAmplitudes [12779] = 8'd131;
   assign soundFileAmplitudes [12780] = 8'd142;
   assign soundFileAmplitudes [12781] = 8'd148;
   assign soundFileAmplitudes [12782] = 8'd111;
   assign soundFileAmplitudes [12783] = 8'd94;
   assign soundFileAmplitudes [12784] = 8'd110;
   assign soundFileAmplitudes [12785] = 8'd114;
   assign soundFileAmplitudes [12786] = 8'd134;
   assign soundFileAmplitudes [12787] = 8'd130;
   assign soundFileAmplitudes [12788] = 8'd126;
   assign soundFileAmplitudes [12789] = 8'd138;
   assign soundFileAmplitudes [12790] = 8'd151;
   assign soundFileAmplitudes [12791] = 8'd153;
   assign soundFileAmplitudes [12792] = 8'd140;
   assign soundFileAmplitudes [12793] = 8'd132;
   assign soundFileAmplitudes [12794] = 8'd123;
   assign soundFileAmplitudes [12795] = 8'd117;
   assign soundFileAmplitudes [12796] = 8'd113;
   assign soundFileAmplitudes [12797] = 8'd103;
   assign soundFileAmplitudes [12798] = 8'd115;
   assign soundFileAmplitudes [12799] = 8'd110;
   assign soundFileAmplitudes [12800] = 8'd114;
   assign soundFileAmplitudes [12801] = 8'd116;
   assign soundFileAmplitudes [12802] = 8'd127;
   assign soundFileAmplitudes [12803] = 8'd143;
   assign soundFileAmplitudes [12804] = 8'd126;
   assign soundFileAmplitudes [12805] = 8'd126;
   assign soundFileAmplitudes [12806] = 8'd115;
   assign soundFileAmplitudes [12807] = 8'd116;
   assign soundFileAmplitudes [12808] = 8'd130;
   assign soundFileAmplitudes [12809] = 8'd147;
   assign soundFileAmplitudes [12810] = 8'd142;
   assign soundFileAmplitudes [12811] = 8'd134;
   assign soundFileAmplitudes [12812] = 8'd133;
   assign soundFileAmplitudes [12813] = 8'd134;
   assign soundFileAmplitudes [12814] = 8'd136;
   assign soundFileAmplitudes [12815] = 8'd137;
   assign soundFileAmplitudes [12816] = 8'd118;
   assign soundFileAmplitudes [12817] = 8'd119;
   assign soundFileAmplitudes [12818] = 8'd121;
   assign soundFileAmplitudes [12819] = 8'd119;
   assign soundFileAmplitudes [12820] = 8'd117;
   assign soundFileAmplitudes [12821] = 8'd93;
   assign soundFileAmplitudes [12822] = 8'd107;
   assign soundFileAmplitudes [12823] = 8'd112;
   assign soundFileAmplitudes [12824] = 8'd126;
   assign soundFileAmplitudes [12825] = 8'd127;
   assign soundFileAmplitudes [12826] = 8'd127;
   assign soundFileAmplitudes [12827] = 8'd124;
   assign soundFileAmplitudes [12828] = 8'd134;
   assign soundFileAmplitudes [12829] = 8'd137;
   assign soundFileAmplitudes [12830] = 8'd132;
   assign soundFileAmplitudes [12831] = 8'd139;
   assign soundFileAmplitudes [12832] = 8'd128;
   assign soundFileAmplitudes [12833] = 8'd116;
   assign soundFileAmplitudes [12834] = 8'd102;
   assign soundFileAmplitudes [12835] = 8'd106;
   assign soundFileAmplitudes [12836] = 8'd132;
   assign soundFileAmplitudes [12837] = 8'd146;
   assign soundFileAmplitudes [12838] = 8'd139;
   assign soundFileAmplitudes [12839] = 8'd128;
   assign soundFileAmplitudes [12840] = 8'd102;
   assign soundFileAmplitudes [12841] = 8'd118;
   assign soundFileAmplitudes [12842] = 8'd127;
   assign soundFileAmplitudes [12843] = 8'd127;
   assign soundFileAmplitudes [12844] = 8'd128;
   assign soundFileAmplitudes [12845] = 8'd130;
   assign soundFileAmplitudes [12846] = 8'd135;
   assign soundFileAmplitudes [12847] = 8'd133;
   assign soundFileAmplitudes [12848] = 8'd130;
   assign soundFileAmplitudes [12849] = 8'd131;
   assign soundFileAmplitudes [12850] = 8'd131;
   assign soundFileAmplitudes [12851] = 8'd127;
   assign soundFileAmplitudes [12852] = 8'd135;
   assign soundFileAmplitudes [12853] = 8'd130;
   assign soundFileAmplitudes [12854] = 8'd126;
   assign soundFileAmplitudes [12855] = 8'd106;
   assign soundFileAmplitudes [12856] = 8'd114;
   assign soundFileAmplitudes [12857] = 8'd131;
   assign soundFileAmplitudes [12858] = 8'd151;
   assign soundFileAmplitudes [12859] = 8'd136;
   assign soundFileAmplitudes [12860] = 8'd108;
   assign soundFileAmplitudes [12861] = 8'd122;
   assign soundFileAmplitudes [12862] = 8'd113;
   assign soundFileAmplitudes [12863] = 8'd112;
   assign soundFileAmplitudes [12864] = 8'd112;
   assign soundFileAmplitudes [12865] = 8'd110;
   assign soundFileAmplitudes [12866] = 8'd114;
   assign soundFileAmplitudes [12867] = 8'd127;
   assign soundFileAmplitudes [12868] = 8'd140;
   assign soundFileAmplitudes [12869] = 8'd148;
   assign soundFileAmplitudes [12870] = 8'd129;
   assign soundFileAmplitudes [12871] = 8'd109;
   assign soundFileAmplitudes [12872] = 8'd124;
   assign soundFileAmplitudes [12873] = 8'd130;
   assign soundFileAmplitudes [12874] = 8'd146;
   assign soundFileAmplitudes [12875] = 8'd137;
   assign soundFileAmplitudes [12876] = 8'd124;
   assign soundFileAmplitudes [12877] = 8'd131;
   assign soundFileAmplitudes [12878] = 8'd119;
   assign soundFileAmplitudes [12879] = 8'd121;
   assign soundFileAmplitudes [12880] = 8'd131;
   assign soundFileAmplitudes [12881] = 8'd129;
   assign soundFileAmplitudes [12882] = 8'd125;
   assign soundFileAmplitudes [12883] = 8'd119;
   assign soundFileAmplitudes [12884] = 8'd117;
   assign soundFileAmplitudes [12885] = 8'd118;
   assign soundFileAmplitudes [12886] = 8'd119;
   assign soundFileAmplitudes [12887] = 8'd129;
   assign soundFileAmplitudes [12888] = 8'd125;
   assign soundFileAmplitudes [12889] = 8'd122;
   assign soundFileAmplitudes [12890] = 8'd118;
   assign soundFileAmplitudes [12891] = 8'd113;
   assign soundFileAmplitudes [12892] = 8'd110;
   assign soundFileAmplitudes [12893] = 8'd125;
   assign soundFileAmplitudes [12894] = 8'd137;
   assign soundFileAmplitudes [12895] = 8'd130;
   assign soundFileAmplitudes [12896] = 8'd143;
   assign soundFileAmplitudes [12897] = 8'd140;
   assign soundFileAmplitudes [12898] = 8'd138;
   assign soundFileAmplitudes [12899] = 8'd126;
   assign soundFileAmplitudes [12900] = 8'd97;
   assign soundFileAmplitudes [12901] = 8'd113;
   assign soundFileAmplitudes [12902] = 8'd133;
   assign soundFileAmplitudes [12903] = 8'd142;
   assign soundFileAmplitudes [12904] = 8'd148;
   assign soundFileAmplitudes [12905] = 8'd135;
   assign soundFileAmplitudes [12906] = 8'd126;
   assign soundFileAmplitudes [12907] = 8'd119;
   assign soundFileAmplitudes [12908] = 8'd126;
   assign soundFileAmplitudes [12909] = 8'd137;
   assign soundFileAmplitudes [12910] = 8'd139;
   assign soundFileAmplitudes [12911] = 8'd134;
   assign soundFileAmplitudes [12912] = 8'd133;
   assign soundFileAmplitudes [12913] = 8'd126;
   assign soundFileAmplitudes [12914] = 8'd117;
   assign soundFileAmplitudes [12915] = 8'd126;
   assign soundFileAmplitudes [12916] = 8'd123;
   assign soundFileAmplitudes [12917] = 8'd117;
   assign soundFileAmplitudes [12918] = 8'd115;
   assign soundFileAmplitudes [12919] = 8'd108;
   assign soundFileAmplitudes [12920] = 8'd108;
   assign soundFileAmplitudes [12921] = 8'd108;
   assign soundFileAmplitudes [12922] = 8'd106;
   assign soundFileAmplitudes [12923] = 8'd111;
   assign soundFileAmplitudes [12924] = 8'd120;
   assign soundFileAmplitudes [12925] = 8'd129;
   assign soundFileAmplitudes [12926] = 8'd136;
   assign soundFileAmplitudes [12927] = 8'd140;
   assign soundFileAmplitudes [12928] = 8'd122;
   assign soundFileAmplitudes [12929] = 8'd118;
   assign soundFileAmplitudes [12930] = 8'd122;
   assign soundFileAmplitudes [12931] = 8'd136;
   assign soundFileAmplitudes [12932] = 8'd143;
   assign soundFileAmplitudes [12933] = 8'd143;
   assign soundFileAmplitudes [12934] = 8'd125;
   assign soundFileAmplitudes [12935] = 8'd119;
   assign soundFileAmplitudes [12936] = 8'd123;
   assign soundFileAmplitudes [12937] = 8'd130;
   assign soundFileAmplitudes [12938] = 8'd156;
   assign soundFileAmplitudes [12939] = 8'd126;
   assign soundFileAmplitudes [12940] = 8'd123;
   assign soundFileAmplitudes [12941] = 8'd131;
   assign soundFileAmplitudes [12942] = 8'd126;
   assign soundFileAmplitudes [12943] = 8'd134;
   assign soundFileAmplitudes [12944] = 8'd132;
   assign soundFileAmplitudes [12945] = 8'd126;
   assign soundFileAmplitudes [12946] = 8'd128;
   assign soundFileAmplitudes [12947] = 8'd120;
   assign soundFileAmplitudes [12948] = 8'd132;
   assign soundFileAmplitudes [12949] = 8'd140;
   assign soundFileAmplitudes [12950] = 8'd122;
   assign soundFileAmplitudes [12951] = 8'd124;
   assign soundFileAmplitudes [12952] = 8'd123;
   assign soundFileAmplitudes [12953] = 8'd124;
   assign soundFileAmplitudes [12954] = 8'd122;
   assign soundFileAmplitudes [12955] = 8'd116;
   assign soundFileAmplitudes [12956] = 8'd116;
   assign soundFileAmplitudes [12957] = 8'd117;
   assign soundFileAmplitudes [12958] = 8'd110;
   assign soundFileAmplitudes [12959] = 8'd113;
   assign soundFileAmplitudes [12960] = 8'd117;
   assign soundFileAmplitudes [12961] = 8'd123;
   assign soundFileAmplitudes [12962] = 8'd131;
   assign soundFileAmplitudes [12963] = 8'd123;
   assign soundFileAmplitudes [12964] = 8'd116;
   assign soundFileAmplitudes [12965] = 8'd115;
   assign soundFileAmplitudes [12966] = 8'd114;
   assign soundFileAmplitudes [12967] = 8'd127;
   assign soundFileAmplitudes [12968] = 8'd134;
   assign soundFileAmplitudes [12969] = 8'd135;
   assign soundFileAmplitudes [12970] = 8'd130;
   assign soundFileAmplitudes [12971] = 8'd120;
   assign soundFileAmplitudes [12972] = 8'd125;
   assign soundFileAmplitudes [12973] = 8'd118;
   assign soundFileAmplitudes [12974] = 8'd120;
   assign soundFileAmplitudes [12975] = 8'd145;
   assign soundFileAmplitudes [12976] = 8'd155;
   assign soundFileAmplitudes [12977] = 8'd167;
   assign soundFileAmplitudes [12978] = 8'd159;
   assign soundFileAmplitudes [12979] = 8'd125;
   assign soundFileAmplitudes [12980] = 8'd125;
   assign soundFileAmplitudes [12981] = 8'd127;
   assign soundFileAmplitudes [12982] = 8'd125;
   assign soundFileAmplitudes [12983] = 8'd117;
   assign soundFileAmplitudes [12984] = 8'd99;
   assign soundFileAmplitudes [12985] = 8'd107;
   assign soundFileAmplitudes [12986] = 8'd110;
   assign soundFileAmplitudes [12987] = 8'd113;
   assign soundFileAmplitudes [12988] = 8'd121;
   assign soundFileAmplitudes [12989] = 8'd123;
   assign soundFileAmplitudes [12990] = 8'd130;
   assign soundFileAmplitudes [12991] = 8'd138;
   assign soundFileAmplitudes [12992] = 8'd133;
   assign soundFileAmplitudes [12993] = 8'd132;
   assign soundFileAmplitudes [12994] = 8'd126;
   assign soundFileAmplitudes [12995] = 8'd114;
   assign soundFileAmplitudes [12996] = 8'd104;
   assign soundFileAmplitudes [12997] = 8'd112;
   assign soundFileAmplitudes [12998] = 8'd115;
   assign soundFileAmplitudes [12999] = 8'd112;
   assign soundFileAmplitudes [13000] = 8'd111;
   assign soundFileAmplitudes [13001] = 8'd111;
   assign soundFileAmplitudes [13002] = 8'd113;
   assign soundFileAmplitudes [13003] = 8'd113;
   assign soundFileAmplitudes [13004] = 8'd132;
   assign soundFileAmplitudes [13005] = 8'd145;
   assign soundFileAmplitudes [13006] = 8'd153;
   assign soundFileAmplitudes [13007] = 8'd142;
   assign soundFileAmplitudes [13008] = 8'd125;
   assign soundFileAmplitudes [13009] = 8'd115;
   assign soundFileAmplitudes [13010] = 8'd123;
   assign soundFileAmplitudes [13011] = 8'd148;
   assign soundFileAmplitudes [13012] = 8'd164;
   assign soundFileAmplitudes [13013] = 8'd148;
   assign soundFileAmplitudes [13014] = 8'd137;
   assign soundFileAmplitudes [13015] = 8'd140;
   assign soundFileAmplitudes [13016] = 8'd164;
   assign soundFileAmplitudes [13017] = 8'd166;
   assign soundFileAmplitudes [13018] = 8'd119;
   assign soundFileAmplitudes [13019] = 8'd102;
   assign soundFileAmplitudes [13020] = 8'd91;
   assign soundFileAmplitudes [13021] = 8'd104;
   assign soundFileAmplitudes [13022] = 8'd113;
   assign soundFileAmplitudes [13023] = 8'd108;
   assign soundFileAmplitudes [13024] = 8'd108;
   assign soundFileAmplitudes [13025] = 8'd114;
   assign soundFileAmplitudes [13026] = 8'd120;
   assign soundFileAmplitudes [13027] = 8'd120;
   assign soundFileAmplitudes [13028] = 8'd116;
   assign soundFileAmplitudes [13029] = 8'd125;
   assign soundFileAmplitudes [13030] = 8'd130;
   assign soundFileAmplitudes [13031] = 8'd127;
   assign soundFileAmplitudes [13032] = 8'd132;
   assign soundFileAmplitudes [13033] = 8'd128;
   assign soundFileAmplitudes [13034] = 8'd129;
   assign soundFileAmplitudes [13035] = 8'd127;
   assign soundFileAmplitudes [13036] = 8'd126;
   assign soundFileAmplitudes [13037] = 8'd123;
   assign soundFileAmplitudes [13038] = 8'd136;
   assign soundFileAmplitudes [13039] = 8'd131;
   assign soundFileAmplitudes [13040] = 8'd121;
   assign soundFileAmplitudes [13041] = 8'd122;
   assign soundFileAmplitudes [13042] = 8'd122;
   assign soundFileAmplitudes [13043] = 8'd125;
   assign soundFileAmplitudes [13044] = 8'd122;
   assign soundFileAmplitudes [13045] = 8'd109;
   assign soundFileAmplitudes [13046] = 8'd110;
   assign soundFileAmplitudes [13047] = 8'd110;
   assign soundFileAmplitudes [13048] = 8'd117;
   assign soundFileAmplitudes [13049] = 8'd137;
   assign soundFileAmplitudes [13050] = 8'd161;
   assign soundFileAmplitudes [13051] = 8'd150;
   assign soundFileAmplitudes [13052] = 8'd137;
   assign soundFileAmplitudes [13053] = 8'd159;
   assign soundFileAmplitudes [13054] = 8'd161;
   assign soundFileAmplitudes [13055] = 8'd167;
   assign soundFileAmplitudes [13056] = 8'd110;
   assign soundFileAmplitudes [13057] = 8'd79;
   assign soundFileAmplitudes [13058] = 8'd103;
   assign soundFileAmplitudes [13059] = 8'd113;
   assign soundFileAmplitudes [13060] = 8'd123;
   assign soundFileAmplitudes [13061] = 8'd117;
   assign soundFileAmplitudes [13062] = 8'd99;
   assign soundFileAmplitudes [13063] = 8'd91;
   assign soundFileAmplitudes [13064] = 8'd99;
   assign soundFileAmplitudes [13065] = 8'd123;
   assign soundFileAmplitudes [13066] = 8'd146;
   assign soundFileAmplitudes [13067] = 8'd140;
   assign soundFileAmplitudes [13068] = 8'd150;
   assign soundFileAmplitudes [13069] = 8'd154;
   assign soundFileAmplitudes [13070] = 8'd142;
   assign soundFileAmplitudes [13071] = 8'd143;
   assign soundFileAmplitudes [13072] = 8'd146;
   assign soundFileAmplitudes [13073] = 8'd139;
   assign soundFileAmplitudes [13074] = 8'd134;
   assign soundFileAmplitudes [13075] = 8'd118;
   assign soundFileAmplitudes [13076] = 8'd103;
   assign soundFileAmplitudes [13077] = 8'd98;
   assign soundFileAmplitudes [13078] = 8'd96;
   assign soundFileAmplitudes [13079] = 8'd99;
   assign soundFileAmplitudes [13080] = 8'd98;
   assign soundFileAmplitudes [13081] = 8'd100;
   assign soundFileAmplitudes [13082] = 8'd97;
   assign soundFileAmplitudes [13083] = 8'd113;
   assign soundFileAmplitudes [13084] = 8'd129;
   assign soundFileAmplitudes [13085] = 8'd138;
   assign soundFileAmplitudes [13086] = 8'd135;
   assign soundFileAmplitudes [13087] = 8'd143;
   assign soundFileAmplitudes [13088] = 8'd170;
   assign soundFileAmplitudes [13089] = 8'd169;
   assign soundFileAmplitudes [13090] = 8'd157;
   assign soundFileAmplitudes [13091] = 8'd166;
   assign soundFileAmplitudes [13092] = 8'd159;
   assign soundFileAmplitudes [13093] = 8'd147;
   assign soundFileAmplitudes [13094] = 8'd115;
   assign soundFileAmplitudes [13095] = 8'd86;
   assign soundFileAmplitudes [13096] = 8'd103;
   assign soundFileAmplitudes [13097] = 8'd107;
   assign soundFileAmplitudes [13098] = 8'd113;
   assign soundFileAmplitudes [13099] = 8'd110;
   assign soundFileAmplitudes [13100] = 8'd102;
   assign soundFileAmplitudes [13101] = 8'd95;
   assign soundFileAmplitudes [13102] = 8'd102;
   assign soundFileAmplitudes [13103] = 8'd118;
   assign soundFileAmplitudes [13104] = 8'd132;
   assign soundFileAmplitudes [13105] = 8'd151;
   assign soundFileAmplitudes [13106] = 8'd159;
   assign soundFileAmplitudes [13107] = 8'd160;
   assign soundFileAmplitudes [13108] = 8'd139;
   assign soundFileAmplitudes [13109] = 8'd116;
   assign soundFileAmplitudes [13110] = 8'd118;
   assign soundFileAmplitudes [13111] = 8'd128;
   assign soundFileAmplitudes [13112] = 8'd124;
   assign soundFileAmplitudes [13113] = 8'd120;
   assign soundFileAmplitudes [13114] = 8'd116;
   assign soundFileAmplitudes [13115] = 8'd111;
   assign soundFileAmplitudes [13116] = 8'd99;
   assign soundFileAmplitudes [13117] = 8'd98;
   assign soundFileAmplitudes [13118] = 8'd94;
   assign soundFileAmplitudes [13119] = 8'd103;
   assign soundFileAmplitudes [13120] = 8'd131;
   assign soundFileAmplitudes [13121] = 8'd140;
   assign soundFileAmplitudes [13122] = 8'd150;
   assign soundFileAmplitudes [13123] = 8'd133;
   assign soundFileAmplitudes [13124] = 8'd122;
   assign soundFileAmplitudes [13125] = 8'd138;
   assign soundFileAmplitudes [13126] = 8'd162;
   assign soundFileAmplitudes [13127] = 8'd170;
   assign soundFileAmplitudes [13128] = 8'd146;
   assign soundFileAmplitudes [13129] = 8'd132;
   assign soundFileAmplitudes [13130] = 8'd124;
   assign soundFileAmplitudes [13131] = 8'd142;
   assign soundFileAmplitudes [13132] = 8'd122;
   assign soundFileAmplitudes [13133] = 8'd87;
   assign soundFileAmplitudes [13134] = 8'd106;
   assign soundFileAmplitudes [13135] = 8'd106;
   assign soundFileAmplitudes [13136] = 8'd110;
   assign soundFileAmplitudes [13137] = 8'd123;
   assign soundFileAmplitudes [13138] = 8'd118;
   assign soundFileAmplitudes [13139] = 8'd110;
   assign soundFileAmplitudes [13140] = 8'd106;
   assign soundFileAmplitudes [13141] = 8'd114;
   assign soundFileAmplitudes [13142] = 8'd132;
   assign soundFileAmplitudes [13143] = 8'd144;
   assign soundFileAmplitudes [13144] = 8'd152;
   assign soundFileAmplitudes [13145] = 8'd161;
   assign soundFileAmplitudes [13146] = 8'd145;
   assign soundFileAmplitudes [13147] = 8'd139;
   assign soundFileAmplitudes [13148] = 8'd139;
   assign soundFileAmplitudes [13149] = 8'd135;
   assign soundFileAmplitudes [13150] = 8'd134;
   assign soundFileAmplitudes [13151] = 8'd123;
   assign soundFileAmplitudes [13152] = 8'd115;
   assign soundFileAmplitudes [13153] = 8'd105;
   assign soundFileAmplitudes [13154] = 8'd87;
   assign soundFileAmplitudes [13155] = 8'd66;
   assign soundFileAmplitudes [13156] = 8'd78;
   assign soundFileAmplitudes [13157] = 8'd105;
   assign soundFileAmplitudes [13158] = 8'd121;
   assign soundFileAmplitudes [13159] = 8'd135;
   assign soundFileAmplitudes [13160] = 8'd140;
   assign soundFileAmplitudes [13161] = 8'd136;
   assign soundFileAmplitudes [13162] = 8'd142;
   assign soundFileAmplitudes [13163] = 8'd138;
   assign soundFileAmplitudes [13164] = 8'd151;
   assign soundFileAmplitudes [13165] = 8'd163;
   assign soundFileAmplitudes [13166] = 8'd147;
   assign soundFileAmplitudes [13167] = 8'd142;
   assign soundFileAmplitudes [13168] = 8'd131;
   assign soundFileAmplitudes [13169] = 8'd145;
   assign soundFileAmplitudes [13170] = 8'd170;
   assign soundFileAmplitudes [13171] = 8'd134;
   assign soundFileAmplitudes [13172] = 8'd101;
   assign soundFileAmplitudes [13173] = 8'd100;
   assign soundFileAmplitudes [13174] = 8'd94;
   assign soundFileAmplitudes [13175] = 8'd106;
   assign soundFileAmplitudes [13176] = 8'd108;
   assign soundFileAmplitudes [13177] = 8'd110;
   assign soundFileAmplitudes [13178] = 8'd109;
   assign soundFileAmplitudes [13179] = 8'd114;
   assign soundFileAmplitudes [13180] = 8'd126;
   assign soundFileAmplitudes [13181] = 8'd127;
   assign soundFileAmplitudes [13182] = 8'd134;
   assign soundFileAmplitudes [13183] = 8'd144;
   assign soundFileAmplitudes [13184] = 8'd148;
   assign soundFileAmplitudes [13185] = 8'd137;
   assign soundFileAmplitudes [13186] = 8'd134;
   assign soundFileAmplitudes [13187] = 8'd128;
   assign soundFileAmplitudes [13188] = 8'd123;
   assign soundFileAmplitudes [13189] = 8'd115;
   assign soundFileAmplitudes [13190] = 8'd105;
   assign soundFileAmplitudes [13191] = 8'd94;
   assign soundFileAmplitudes [13192] = 8'd97;
   assign soundFileAmplitudes [13193] = 8'd102;
   assign soundFileAmplitudes [13194] = 8'd103;
   assign soundFileAmplitudes [13195] = 8'd113;
   assign soundFileAmplitudes [13196] = 8'd112;
   assign soundFileAmplitudes [13197] = 8'd122;
   assign soundFileAmplitudes [13198] = 8'd142;
   assign soundFileAmplitudes [13199] = 8'd162;
   assign soundFileAmplitudes [13200] = 8'd163;
   assign soundFileAmplitudes [13201] = 8'd154;
   assign soundFileAmplitudes [13202] = 8'd148;
   assign soundFileAmplitudes [13203] = 8'd165;
   assign soundFileAmplitudes [13204] = 8'd154;
   assign soundFileAmplitudes [13205] = 8'd147;
   assign soundFileAmplitudes [13206] = 8'd146;
   assign soundFileAmplitudes [13207] = 8'd153;
   assign soundFileAmplitudes [13208] = 8'd164;
   assign soundFileAmplitudes [13209] = 8'd120;
   assign soundFileAmplitudes [13210] = 8'd92;
   assign soundFileAmplitudes [13211] = 8'd82;
   assign soundFileAmplitudes [13212] = 8'd82;
   assign soundFileAmplitudes [13213] = 8'd92;
   assign soundFileAmplitudes [13214] = 8'd102;
   assign soundFileAmplitudes [13215] = 8'd103;
   assign soundFileAmplitudes [13216] = 8'd110;
   assign soundFileAmplitudes [13217] = 8'd105;
   assign soundFileAmplitudes [13218] = 8'd108;
   assign soundFileAmplitudes [13219] = 8'd124;
   assign soundFileAmplitudes [13220] = 8'd134;
   assign soundFileAmplitudes [13221] = 8'd143;
   assign soundFileAmplitudes [13222] = 8'd153;
   assign soundFileAmplitudes [13223] = 8'd150;
   assign soundFileAmplitudes [13224] = 8'd140;
   assign soundFileAmplitudes [13225] = 8'd137;
   assign soundFileAmplitudes [13226] = 8'd131;
   assign soundFileAmplitudes [13227] = 8'd116;
   assign soundFileAmplitudes [13228] = 8'd88;
   assign soundFileAmplitudes [13229] = 8'd91;
   assign soundFileAmplitudes [13230] = 8'd101;
   assign soundFileAmplitudes [13231] = 8'd110;
   assign soundFileAmplitudes [13232] = 8'd115;
   assign soundFileAmplitudes [13233] = 8'd115;
   assign soundFileAmplitudes [13234] = 8'd132;
   assign soundFileAmplitudes [13235] = 8'd150;
   assign soundFileAmplitudes [13236] = 8'd165;
   assign soundFileAmplitudes [13237] = 8'd164;
   assign soundFileAmplitudes [13238] = 8'd148;
   assign soundFileAmplitudes [13239] = 8'd151;
   assign soundFileAmplitudes [13240] = 8'd143;
   assign soundFileAmplitudes [13241] = 8'd148;
   assign soundFileAmplitudes [13242] = 8'd163;
   assign soundFileAmplitudes [13243] = 8'd165;
   assign soundFileAmplitudes [13244] = 8'd154;
   assign soundFileAmplitudes [13245] = 8'd134;
   assign soundFileAmplitudes [13246] = 8'd127;
   assign soundFileAmplitudes [13247] = 8'd129;
   assign soundFileAmplitudes [13248] = 8'd102;
   assign soundFileAmplitudes [13249] = 8'd65;
   assign soundFileAmplitudes [13250] = 8'd70;
   assign soundFileAmplitudes [13251] = 8'd79;
   assign soundFileAmplitudes [13252] = 8'd93;
   assign soundFileAmplitudes [13253] = 8'd98;
   assign soundFileAmplitudes [13254] = 8'd83;
   assign soundFileAmplitudes [13255] = 8'd80;
   assign soundFileAmplitudes [13256] = 8'd93;
   assign soundFileAmplitudes [13257] = 8'd107;
   assign soundFileAmplitudes [13258] = 8'd132;
   assign soundFileAmplitudes [13259] = 8'd142;
   assign soundFileAmplitudes [13260] = 8'd153;
   assign soundFileAmplitudes [13261] = 8'd160;
   assign soundFileAmplitudes [13262] = 8'd152;
   assign soundFileAmplitudes [13263] = 8'd133;
   assign soundFileAmplitudes [13264] = 8'd117;
   assign soundFileAmplitudes [13265] = 8'd133;
   assign soundFileAmplitudes [13266] = 8'd141;
   assign soundFileAmplitudes [13267] = 8'd132;
   assign soundFileAmplitudes [13268] = 8'd133;
   assign soundFileAmplitudes [13269] = 8'd126;
   assign soundFileAmplitudes [13270] = 8'd127;
   assign soundFileAmplitudes [13271] = 8'd144;
   assign soundFileAmplitudes [13272] = 8'd147;
   assign soundFileAmplitudes [13273] = 8'd158;
   assign soundFileAmplitudes [13274] = 8'd145;
   assign soundFileAmplitudes [13275] = 8'd142;
   assign soundFileAmplitudes [13276] = 8'd144;
   assign soundFileAmplitudes [13277] = 8'd138;
   assign soundFileAmplitudes [13278] = 8'd142;
   assign soundFileAmplitudes [13279] = 8'd135;
   assign soundFileAmplitudes [13280] = 8'd134;
   assign soundFileAmplitudes [13281] = 8'd131;
   assign soundFileAmplitudes [13282] = 8'd122;
   assign soundFileAmplitudes [13283] = 8'd127;
   assign soundFileAmplitudes [13284] = 8'd114;
   assign soundFileAmplitudes [13285] = 8'd113;
   assign soundFileAmplitudes [13286] = 8'd109;
   assign soundFileAmplitudes [13287] = 8'd87;
   assign soundFileAmplitudes [13288] = 8'd100;
   assign soundFileAmplitudes [13289] = 8'd85;
   assign soundFileAmplitudes [13290] = 8'd68;
   assign soundFileAmplitudes [13291] = 8'd71;
   assign soundFileAmplitudes [13292] = 8'd81;
   assign soundFileAmplitudes [13293] = 8'd91;
   assign soundFileAmplitudes [13294] = 8'd113;
   assign soundFileAmplitudes [13295] = 8'd124;
   assign soundFileAmplitudes [13296] = 8'd124;
   assign soundFileAmplitudes [13297] = 8'd135;
   assign soundFileAmplitudes [13298] = 8'd145;
   assign soundFileAmplitudes [13299] = 8'd153;
   assign soundFileAmplitudes [13300] = 8'd168;
   assign soundFileAmplitudes [13301] = 8'd178;
   assign soundFileAmplitudes [13302] = 8'd163;
   assign soundFileAmplitudes [13303] = 8'd158;
   assign soundFileAmplitudes [13304] = 8'd152;
   assign soundFileAmplitudes [13305] = 8'd146;
   assign soundFileAmplitudes [13306] = 8'd145;
   assign soundFileAmplitudes [13307] = 8'd153;
   assign soundFileAmplitudes [13308] = 8'd143;
   assign soundFileAmplitudes [13309] = 8'd131;
   assign soundFileAmplitudes [13310] = 8'd112;
   assign soundFileAmplitudes [13311] = 8'd101;
   assign soundFileAmplitudes [13312] = 8'd105;
   assign soundFileAmplitudes [13313] = 8'd109;
   assign soundFileAmplitudes [13314] = 8'd122;
   assign soundFileAmplitudes [13315] = 8'd135;
   assign soundFileAmplitudes [13316] = 8'd142;
   assign soundFileAmplitudes [13317] = 8'd141;
   assign soundFileAmplitudes [13318] = 8'd148;
   assign soundFileAmplitudes [13319] = 8'd148;
   assign soundFileAmplitudes [13320] = 8'd142;
   assign soundFileAmplitudes [13321] = 8'd115;
   assign soundFileAmplitudes [13322] = 8'd116;
   assign soundFileAmplitudes [13323] = 8'd122;
   assign soundFileAmplitudes [13324] = 8'd116;
   assign soundFileAmplitudes [13325] = 8'd102;
   assign soundFileAmplitudes [13326] = 8'd62;
   assign soundFileAmplitudes [13327] = 8'd61;
   assign soundFileAmplitudes [13328] = 8'd80;
   assign soundFileAmplitudes [13329] = 8'd81;
   assign soundFileAmplitudes [13330] = 8'd71;
   assign soundFileAmplitudes [13331] = 8'd59;
   assign soundFileAmplitudes [13332] = 8'd68;
   assign soundFileAmplitudes [13333] = 8'd92;
   assign soundFileAmplitudes [13334] = 8'd107;
   assign soundFileAmplitudes [13335] = 8'd126;
   assign soundFileAmplitudes [13336] = 8'd143;
   assign soundFileAmplitudes [13337] = 8'd170;
   assign soundFileAmplitudes [13338] = 8'd181;
   assign soundFileAmplitudes [13339] = 8'd204;
   assign soundFileAmplitudes [13340] = 8'd219;
   assign soundFileAmplitudes [13341] = 8'd196;
   assign soundFileAmplitudes [13342] = 8'd181;
   assign soundFileAmplitudes [13343] = 8'd175;
   assign soundFileAmplitudes [13344] = 8'd175;
   assign soundFileAmplitudes [13345] = 8'd167;
   assign soundFileAmplitudes [13346] = 8'd146;
   assign soundFileAmplitudes [13347] = 8'd131;
   assign soundFileAmplitudes [13348] = 8'd124;
   assign soundFileAmplitudes [13349] = 8'd112;
   assign soundFileAmplitudes [13350] = 8'd107;
   assign soundFileAmplitudes [13351] = 8'd104;
   assign soundFileAmplitudes [13352] = 8'd107;
   assign soundFileAmplitudes [13353] = 8'd112;
   assign soundFileAmplitudes [13354] = 8'd108;
   assign soundFileAmplitudes [13355] = 8'd113;
   assign soundFileAmplitudes [13356] = 8'd116;
   assign soundFileAmplitudes [13357] = 8'd114;
   assign soundFileAmplitudes [13358] = 8'd111;
   assign soundFileAmplitudes [13359] = 8'd125;
   assign soundFileAmplitudes [13360] = 8'd128;
   assign soundFileAmplitudes [13361] = 8'd109;
   assign soundFileAmplitudes [13362] = 8'd104;
   assign soundFileAmplitudes [13363] = 8'd88;
   assign soundFileAmplitudes [13364] = 8'd100;
   assign soundFileAmplitudes [13365] = 8'd98;
   assign soundFileAmplitudes [13366] = 8'd67;
   assign soundFileAmplitudes [13367] = 8'd80;
   assign soundFileAmplitudes [13368] = 8'd101;
   assign soundFileAmplitudes [13369] = 8'd105;
   assign soundFileAmplitudes [13370] = 8'd89;
   assign soundFileAmplitudes [13371] = 8'd79;
   assign soundFileAmplitudes [13372] = 8'd95;
   assign soundFileAmplitudes [13373] = 8'd118;
   assign soundFileAmplitudes [13374] = 8'd156;
   assign soundFileAmplitudes [13375] = 8'd164;
   assign soundFileAmplitudes [13376] = 8'd170;
   assign soundFileAmplitudes [13377] = 8'd181;
   assign soundFileAmplitudes [13378] = 8'd190;
   assign soundFileAmplitudes [13379] = 8'd204;
   assign soundFileAmplitudes [13380] = 8'd213;
   assign soundFileAmplitudes [13381] = 8'd213;
   assign soundFileAmplitudes [13382] = 8'd175;
   assign soundFileAmplitudes [13383] = 8'd157;
   assign soundFileAmplitudes [13384] = 8'd133;
   assign soundFileAmplitudes [13385] = 8'd127;
   assign soundFileAmplitudes [13386] = 8'd124;
   assign soundFileAmplitudes [13387] = 8'd117;
   assign soundFileAmplitudes [13388] = 8'd106;
   assign soundFileAmplitudes [13389] = 8'd88;
   assign soundFileAmplitudes [13390] = 8'd95;
   assign soundFileAmplitudes [13391] = 8'd87;
   assign soundFileAmplitudes [13392] = 8'd93;
   assign soundFileAmplitudes [13393] = 8'd106;
   assign soundFileAmplitudes [13394] = 8'd112;
   assign soundFileAmplitudes [13395] = 8'd118;
   assign soundFileAmplitudes [13396] = 8'd124;
   assign soundFileAmplitudes [13397] = 8'd120;
   assign soundFileAmplitudes [13398] = 8'd121;
   assign soundFileAmplitudes [13399] = 8'd115;
   assign soundFileAmplitudes [13400] = 8'd117;
   assign soundFileAmplitudes [13401] = 8'd106;
   assign soundFileAmplitudes [13402] = 8'd105;
   assign soundFileAmplitudes [13403] = 8'd111;
   assign soundFileAmplitudes [13404] = 8'd110;
   assign soundFileAmplitudes [13405] = 8'd116;
   assign soundFileAmplitudes [13406] = 8'd104;
   assign soundFileAmplitudes [13407] = 8'd108;
   assign soundFileAmplitudes [13408] = 8'd104;
   assign soundFileAmplitudes [13409] = 8'd104;
   assign soundFileAmplitudes [13410] = 8'd94;
   assign soundFileAmplitudes [13411] = 8'd86;
   assign soundFileAmplitudes [13412] = 8'd96;
   assign soundFileAmplitudes [13413] = 8'd116;
   assign soundFileAmplitudes [13414] = 8'd139;
   assign soundFileAmplitudes [13415] = 8'd140;
   assign soundFileAmplitudes [13416] = 8'd157;
   assign soundFileAmplitudes [13417] = 8'd168;
   assign soundFileAmplitudes [13418] = 8'd189;
   assign soundFileAmplitudes [13419] = 8'd203;
   assign soundFileAmplitudes [13420] = 8'd200;
   assign soundFileAmplitudes [13421] = 8'd194;
   assign soundFileAmplitudes [13422] = 8'd166;
   assign soundFileAmplitudes [13423] = 8'd150;
   assign soundFileAmplitudes [13424] = 8'd139;
   assign soundFileAmplitudes [13425] = 8'd140;
   assign soundFileAmplitudes [13426] = 8'd133;
   assign soundFileAmplitudes [13427] = 8'd120;
   assign soundFileAmplitudes [13428] = 8'd109;
   assign soundFileAmplitudes [13429] = 8'd97;
   assign soundFileAmplitudes [13430] = 8'd93;
   assign soundFileAmplitudes [13431] = 8'd84;
   assign soundFileAmplitudes [13432] = 8'd77;
   assign soundFileAmplitudes [13433] = 8'd76;
   assign soundFileAmplitudes [13434] = 8'd89;
   assign soundFileAmplitudes [13435] = 8'd102;
   assign soundFileAmplitudes [13436] = 8'd121;
   assign soundFileAmplitudes [13437] = 8'd141;
   assign soundFileAmplitudes [13438] = 8'd141;
   assign soundFileAmplitudes [13439] = 8'd135;
   assign soundFileAmplitudes [13440] = 8'd135;
   assign soundFileAmplitudes [13441] = 8'd128;
   assign soundFileAmplitudes [13442] = 8'd125;
   assign soundFileAmplitudes [13443] = 8'd129;
   assign soundFileAmplitudes [13444] = 8'd132;
   assign soundFileAmplitudes [13445] = 8'd138;
   assign soundFileAmplitudes [13446] = 8'd116;
   assign soundFileAmplitudes [13447] = 8'd96;
   assign soundFileAmplitudes [13448] = 8'd105;
   assign soundFileAmplitudes [13449] = 8'd115;
   assign soundFileAmplitudes [13450] = 8'd114;
   assign soundFileAmplitudes [13451] = 8'd106;
   assign soundFileAmplitudes [13452] = 8'd87;
   assign soundFileAmplitudes [13453] = 8'd85;
   assign soundFileAmplitudes [13454] = 8'd97;
   assign soundFileAmplitudes [13455] = 8'd123;
   assign soundFileAmplitudes [13456] = 8'd157;
   assign soundFileAmplitudes [13457] = 8'd168;
   assign soundFileAmplitudes [13458] = 8'd185;
   assign soundFileAmplitudes [13459] = 8'd182;
   assign soundFileAmplitudes [13460] = 8'd181;
   assign soundFileAmplitudes [13461] = 8'd174;
   assign soundFileAmplitudes [13462] = 8'd158;
   assign soundFileAmplitudes [13463] = 8'd154;
   assign soundFileAmplitudes [13464] = 8'd149;
   assign soundFileAmplitudes [13465] = 8'd138;
   assign soundFileAmplitudes [13466] = 8'd129;
   assign soundFileAmplitudes [13467] = 8'd112;
   assign soundFileAmplitudes [13468] = 8'd89;
   assign soundFileAmplitudes [13469] = 8'd78;
   assign soundFileAmplitudes [13470] = 8'd74;
   assign soundFileAmplitudes [13471] = 8'd87;
   assign soundFileAmplitudes [13472] = 8'd93;
   assign soundFileAmplitudes [13473] = 8'd103;
   assign soundFileAmplitudes [13474] = 8'd112;
   assign soundFileAmplitudes [13475] = 8'd120;
   assign soundFileAmplitudes [13476] = 8'd135;
   assign soundFileAmplitudes [13477] = 8'd140;
   assign soundFileAmplitudes [13478] = 8'd137;
   assign soundFileAmplitudes [13479] = 8'd141;
   assign soundFileAmplitudes [13480] = 8'd140;
   assign soundFileAmplitudes [13481] = 8'd138;
   assign soundFileAmplitudes [13482] = 8'd129;
   assign soundFileAmplitudes [13483] = 8'd125;
   assign soundFileAmplitudes [13484] = 8'd124;
   assign soundFileAmplitudes [13485] = 8'd123;
   assign soundFileAmplitudes [13486] = 8'd119;
   assign soundFileAmplitudes [13487] = 8'd113;
   assign soundFileAmplitudes [13488] = 8'd107;
   assign soundFileAmplitudes [13489] = 8'd102;
   assign soundFileAmplitudes [13490] = 8'd111;
   assign soundFileAmplitudes [13491] = 8'd117;
   assign soundFileAmplitudes [13492] = 8'd122;
   assign soundFileAmplitudes [13493] = 8'd127;
   assign soundFileAmplitudes [13494] = 8'd120;
   assign soundFileAmplitudes [13495] = 8'd112;
   assign soundFileAmplitudes [13496] = 8'd129;
   assign soundFileAmplitudes [13497] = 8'd133;
   assign soundFileAmplitudes [13498] = 8'd154;
   assign soundFileAmplitudes [13499] = 8'd163;
   assign soundFileAmplitudes [13500] = 8'd154;
   assign soundFileAmplitudes [13501] = 8'd154;
   assign soundFileAmplitudes [13502] = 8'd142;
   assign soundFileAmplitudes [13503] = 8'd143;
   assign soundFileAmplitudes [13504] = 8'd131;
   assign soundFileAmplitudes [13505] = 8'd119;
   assign soundFileAmplitudes [13506] = 8'd116;
   assign soundFileAmplitudes [13507] = 8'd106;
   assign soundFileAmplitudes [13508] = 8'd109;
   assign soundFileAmplitudes [13509] = 8'd116;
   assign soundFileAmplitudes [13510] = 8'd120;
   assign soundFileAmplitudes [13511] = 8'd126;
   assign soundFileAmplitudes [13512] = 8'd129;
   assign soundFileAmplitudes [13513] = 8'd126;
   assign soundFileAmplitudes [13514] = 8'd121;
   assign soundFileAmplitudes [13515] = 8'd128;
   assign soundFileAmplitudes [13516] = 8'd130;
   assign soundFileAmplitudes [13517] = 8'd132;
   assign soundFileAmplitudes [13518] = 8'd136;
   assign soundFileAmplitudes [13519] = 8'd146;
   assign soundFileAmplitudes [13520] = 8'd145;
   assign soundFileAmplitudes [13521] = 8'd134;
   assign soundFileAmplitudes [13522] = 8'd123;
   assign soundFileAmplitudes [13523] = 8'd119;
   assign soundFileAmplitudes [13524] = 8'd123;
   assign soundFileAmplitudes [13525] = 8'd119;
   assign soundFileAmplitudes [13526] = 8'd110;
   assign soundFileAmplitudes [13527] = 8'd107;
   assign soundFileAmplitudes [13528] = 8'd116;
   assign soundFileAmplitudes [13529] = 8'd129;
   assign soundFileAmplitudes [13530] = 8'd128;
   assign soundFileAmplitudes [13531] = 8'd129;
   assign soundFileAmplitudes [13532] = 8'd121;
   assign soundFileAmplitudes [13533] = 8'd106;
   assign soundFileAmplitudes [13534] = 8'd109;
   assign soundFileAmplitudes [13535] = 8'd97;
   assign soundFileAmplitudes [13536] = 8'd107;
   assign soundFileAmplitudes [13537] = 8'd115;
   assign soundFileAmplitudes [13538] = 8'd115;
   assign soundFileAmplitudes [13539] = 8'd119;
   assign soundFileAmplitudes [13540] = 8'd116;
   assign soundFileAmplitudes [13541] = 8'd117;
   assign soundFileAmplitudes [13542] = 8'd118;
   assign soundFileAmplitudes [13543] = 8'd130;
   assign soundFileAmplitudes [13544] = 8'd140;
   assign soundFileAmplitudes [13545] = 8'd139;
   assign soundFileAmplitudes [13546] = 8'd140;
   assign soundFileAmplitudes [13547] = 8'd135;
   assign soundFileAmplitudes [13548] = 8'd123;
   assign soundFileAmplitudes [13549] = 8'd120;
   assign soundFileAmplitudes [13550] = 8'd121;
   assign soundFileAmplitudes [13551] = 8'd126;
   assign soundFileAmplitudes [13552] = 8'd133;
   assign soundFileAmplitudes [13553] = 8'd139;
   assign soundFileAmplitudes [13554] = 8'd145;
   assign soundFileAmplitudes [13555] = 8'd150;
   assign soundFileAmplitudes [13556] = 8'd143;
   assign soundFileAmplitudes [13557] = 8'd137;
   assign soundFileAmplitudes [13558] = 8'd126;
   assign soundFileAmplitudes [13559] = 8'd123;
   assign soundFileAmplitudes [13560] = 8'd120;
   assign soundFileAmplitudes [13561] = 8'd131;
   assign soundFileAmplitudes [13562] = 8'd147;
   assign soundFileAmplitudes [13563] = 8'd149;
   assign soundFileAmplitudes [13564] = 8'd154;
   assign soundFileAmplitudes [13565] = 8'd137;
   assign soundFileAmplitudes [13566] = 8'd117;
   assign soundFileAmplitudes [13567] = 8'd104;
   assign soundFileAmplitudes [13568] = 8'd104;
   assign soundFileAmplitudes [13569] = 8'd119;
   assign soundFileAmplitudes [13570] = 8'd120;
   assign soundFileAmplitudes [13571] = 8'd117;
   assign soundFileAmplitudes [13572] = 8'd116;
   assign soundFileAmplitudes [13573] = 8'd97;
   assign soundFileAmplitudes [13574] = 8'd94;
   assign soundFileAmplitudes [13575] = 8'd88;
   assign soundFileAmplitudes [13576] = 8'd98;
   assign soundFileAmplitudes [13577] = 8'd117;
   assign soundFileAmplitudes [13578] = 8'd133;
   assign soundFileAmplitudes [13579] = 8'd143;
   assign soundFileAmplitudes [13580] = 8'd120;
   assign soundFileAmplitudes [13581] = 8'd108;
   assign soundFileAmplitudes [13582] = 8'd107;
   assign soundFileAmplitudes [13583] = 8'd114;
   assign soundFileAmplitudes [13584] = 8'd120;
   assign soundFileAmplitudes [13585] = 8'd132;
   assign soundFileAmplitudes [13586] = 8'd141;
   assign soundFileAmplitudes [13587] = 8'd146;
   assign soundFileAmplitudes [13588] = 8'd146;
   assign soundFileAmplitudes [13589] = 8'd149;
   assign soundFileAmplitudes [13590] = 8'd154;
   assign soundFileAmplitudes [13591] = 8'd142;
   assign soundFileAmplitudes [13592] = 8'd139;
   assign soundFileAmplitudes [13593] = 8'd142;
   assign soundFileAmplitudes [13594] = 8'd153;
   assign soundFileAmplitudes [13595] = 8'd149;
   assign soundFileAmplitudes [13596] = 8'd149;
   assign soundFileAmplitudes [13597] = 8'd152;
   assign soundFileAmplitudes [13598] = 8'd139;
   assign soundFileAmplitudes [13599] = 8'd136;
   assign soundFileAmplitudes [13600] = 8'd126;
   assign soundFileAmplitudes [13601] = 8'd128;
   assign soundFileAmplitudes [13602] = 8'd138;
   assign soundFileAmplitudes [13603] = 8'd132;
   assign soundFileAmplitudes [13604] = 8'd123;
   assign soundFileAmplitudes [13605] = 8'd113;
   assign soundFileAmplitudes [13606] = 8'd106;
   assign soundFileAmplitudes [13607] = 8'd125;
   assign soundFileAmplitudes [13608] = 8'd119;
   assign soundFileAmplitudes [13609] = 8'd103;
   assign soundFileAmplitudes [13610] = 8'd103;
   assign soundFileAmplitudes [13611] = 8'd89;
   assign soundFileAmplitudes [13612] = 8'd95;
   assign soundFileAmplitudes [13613] = 8'd96;
   assign soundFileAmplitudes [13614] = 8'd97;
   assign soundFileAmplitudes [13615] = 8'd98;
   assign soundFileAmplitudes [13616] = 8'd103;
   assign soundFileAmplitudes [13617] = 8'd111;
   assign soundFileAmplitudes [13618] = 8'd104;
   assign soundFileAmplitudes [13619] = 8'd101;
   assign soundFileAmplitudes [13620] = 8'd99;
   assign soundFileAmplitudes [13621] = 8'd99;
   assign soundFileAmplitudes [13622] = 8'd117;
   assign soundFileAmplitudes [13623] = 8'd133;
   assign soundFileAmplitudes [13624] = 8'd138;
   assign soundFileAmplitudes [13625] = 8'd157;
   assign soundFileAmplitudes [13626] = 8'd169;
   assign soundFileAmplitudes [13627] = 8'd168;
   assign soundFileAmplitudes [13628] = 8'd169;
   assign soundFileAmplitudes [13629] = 8'd153;
   assign soundFileAmplitudes [13630] = 8'd137;
   assign soundFileAmplitudes [13631] = 8'd139;
   assign soundFileAmplitudes [13632] = 8'd155;
   assign soundFileAmplitudes [13633] = 8'd166;
   assign soundFileAmplitudes [13634] = 8'd162;
   assign soundFileAmplitudes [13635] = 8'd145;
   assign soundFileAmplitudes [13636] = 8'd129;
   assign soundFileAmplitudes [13637] = 8'd132;
   assign soundFileAmplitudes [13638] = 8'd128;
   assign soundFileAmplitudes [13639] = 8'd135;
   assign soundFileAmplitudes [13640] = 8'd122;
   assign soundFileAmplitudes [13641] = 8'd121;
   assign soundFileAmplitudes [13642] = 8'd132;
   assign soundFileAmplitudes [13643] = 8'd123;
   assign soundFileAmplitudes [13644] = 8'd107;
   assign soundFileAmplitudes [13645] = 8'd102;
   assign soundFileAmplitudes [13646] = 8'd98;
   assign soundFileAmplitudes [13647] = 8'd109;
   assign soundFileAmplitudes [13648] = 8'd122;
   assign soundFileAmplitudes [13649] = 8'd112;
   assign soundFileAmplitudes [13650] = 8'd111;
   assign soundFileAmplitudes [13651] = 8'd99;
   assign soundFileAmplitudes [13652] = 8'd90;
   assign soundFileAmplitudes [13653] = 8'd80;
   assign soundFileAmplitudes [13654] = 8'd80;
   assign soundFileAmplitudes [13655] = 8'd102;
   assign soundFileAmplitudes [13656] = 8'd113;
   assign soundFileAmplitudes [13657] = 8'd115;
   assign soundFileAmplitudes [13658] = 8'd120;
   assign soundFileAmplitudes [13659] = 8'd118;
   assign soundFileAmplitudes [13660] = 8'd129;
   assign soundFileAmplitudes [13661] = 8'd144;
   assign soundFileAmplitudes [13662] = 8'd157;
   assign soundFileAmplitudes [13663] = 8'd156;
   assign soundFileAmplitudes [13664] = 8'd154;
   assign soundFileAmplitudes [13665] = 8'd148;
   assign soundFileAmplitudes [13666] = 8'd149;
   assign soundFileAmplitudes [13667] = 8'd161;
   assign soundFileAmplitudes [13668] = 8'd150;
   assign soundFileAmplitudes [13669] = 8'd139;
   assign soundFileAmplitudes [13670] = 8'd126;
   assign soundFileAmplitudes [13671] = 8'd117;
   assign soundFileAmplitudes [13672] = 8'd119;
   assign soundFileAmplitudes [13673] = 8'd116;
   assign soundFileAmplitudes [13674] = 8'd118;
   assign soundFileAmplitudes [13675] = 8'd123;
   assign soundFileAmplitudes [13676] = 8'd126;
   assign soundFileAmplitudes [13677] = 8'd141;
   assign soundFileAmplitudes [13678] = 8'd138;
   assign soundFileAmplitudes [13679] = 8'd130;
   assign soundFileAmplitudes [13680] = 8'd116;
   assign soundFileAmplitudes [13681] = 8'd118;
   assign soundFileAmplitudes [13682] = 8'd137;
   assign soundFileAmplitudes [13683] = 8'd152;
   assign soundFileAmplitudes [13684] = 8'd150;
   assign soundFileAmplitudes [13685] = 8'd137;
   assign soundFileAmplitudes [13686] = 8'd115;
   assign soundFileAmplitudes [13687] = 8'd120;
   assign soundFileAmplitudes [13688] = 8'd129;
   assign soundFileAmplitudes [13689] = 8'd110;
   assign soundFileAmplitudes [13690] = 8'd111;
   assign soundFileAmplitudes [13691] = 8'd109;
   assign soundFileAmplitudes [13692] = 8'd118;
   assign soundFileAmplitudes [13693] = 8'd110;
   assign soundFileAmplitudes [13694] = 8'd114;
   assign soundFileAmplitudes [13695] = 8'd120;
   assign soundFileAmplitudes [13696] = 8'd122;
   assign soundFileAmplitudes [13697] = 8'd120;
   assign soundFileAmplitudes [13698] = 8'd99;
   assign soundFileAmplitudes [13699] = 8'd97;
   assign soundFileAmplitudes [13700] = 8'd108;
   assign soundFileAmplitudes [13701] = 8'd109;
   assign soundFileAmplitudes [13702] = 8'd114;
   assign soundFileAmplitudes [13703] = 8'd132;
   assign soundFileAmplitudes [13704] = 8'd131;
   assign soundFileAmplitudes [13705] = 8'd132;
   assign soundFileAmplitudes [13706] = 8'd136;
   assign soundFileAmplitudes [13707] = 8'd142;
   assign soundFileAmplitudes [13708] = 8'd136;
   assign soundFileAmplitudes [13709] = 8'd117;
   assign soundFileAmplitudes [13710] = 8'd103;
   assign soundFileAmplitudes [13711] = 8'd110;
   assign soundFileAmplitudes [13712] = 8'd124;
   assign soundFileAmplitudes [13713] = 8'd141;
   assign soundFileAmplitudes [13714] = 8'd141;
   assign soundFileAmplitudes [13715] = 8'd127;
   assign soundFileAmplitudes [13716] = 8'd130;
   assign soundFileAmplitudes [13717] = 8'd126;
   assign soundFileAmplitudes [13718] = 8'd124;
   assign soundFileAmplitudes [13719] = 8'd137;
   assign soundFileAmplitudes [13720] = 8'd160;
   assign soundFileAmplitudes [13721] = 8'd156;
   assign soundFileAmplitudes [13722] = 8'd151;
   assign soundFileAmplitudes [13723] = 8'd145;
   assign soundFileAmplitudes [13724] = 8'd136;
   assign soundFileAmplitudes [13725] = 8'd137;
   assign soundFileAmplitudes [13726] = 8'd130;
   assign soundFileAmplitudes [13727] = 8'd122;
   assign soundFileAmplitudes [13728] = 8'd135;
   assign soundFileAmplitudes [13729] = 8'd135;
   assign soundFileAmplitudes [13730] = 8'd134;
   assign soundFileAmplitudes [13731] = 8'd143;
   assign soundFileAmplitudes [13732] = 8'd131;
   assign soundFileAmplitudes [13733] = 8'd124;
   assign soundFileAmplitudes [13734] = 8'd94;
   assign soundFileAmplitudes [13735] = 8'd78;
   assign soundFileAmplitudes [13736] = 8'd84;
   assign soundFileAmplitudes [13737] = 8'd98;
   assign soundFileAmplitudes [13738] = 8'd115;
   assign soundFileAmplitudes [13739] = 8'd125;
   assign soundFileAmplitudes [13740] = 8'd127;
   assign soundFileAmplitudes [13741] = 8'd135;
   assign soundFileAmplitudes [13742] = 8'd134;
   assign soundFileAmplitudes [13743] = 8'd140;
   assign soundFileAmplitudes [13744] = 8'd143;
   assign soundFileAmplitudes [13745] = 8'd132;
   assign soundFileAmplitudes [13746] = 8'd123;
   assign soundFileAmplitudes [13747] = 8'd114;
   assign soundFileAmplitudes [13748] = 8'd117;
   assign soundFileAmplitudes [13749] = 8'd118;
   assign soundFileAmplitudes [13750] = 8'd107;
   assign soundFileAmplitudes [13751] = 8'd107;
   assign soundFileAmplitudes [13752] = 8'd109;
   assign soundFileAmplitudes [13753] = 8'd112;
   assign soundFileAmplitudes [13754] = 8'd120;
   assign soundFileAmplitudes [13755] = 8'd124;
   assign soundFileAmplitudes [13756] = 8'd127;
   assign soundFileAmplitudes [13757] = 8'd126;
   assign soundFileAmplitudes [13758] = 8'd140;
   assign soundFileAmplitudes [13759] = 8'd140;
   assign soundFileAmplitudes [13760] = 8'd151;
   assign soundFileAmplitudes [13761] = 8'd152;
   assign soundFileAmplitudes [13762] = 8'd152;
   assign soundFileAmplitudes [13763] = 8'd146;
   assign soundFileAmplitudes [13764] = 8'd124;
   assign soundFileAmplitudes [13765] = 8'd120;
   assign soundFileAmplitudes [13766] = 8'd145;
   assign soundFileAmplitudes [13767] = 8'd139;
   assign soundFileAmplitudes [13768] = 8'd113;
   assign soundFileAmplitudes [13769] = 8'd128;
   assign soundFileAmplitudes [13770] = 8'd123;
   assign soundFileAmplitudes [13771] = 8'd123;
   assign soundFileAmplitudes [13772] = 8'd100;
   assign soundFileAmplitudes [13773] = 8'd86;
   assign soundFileAmplitudes [13774] = 8'd99;
   assign soundFileAmplitudes [13775] = 8'd116;
   assign soundFileAmplitudes [13776] = 8'd132;
   assign soundFileAmplitudes [13777] = 8'd128;
   assign soundFileAmplitudes [13778] = 8'd125;
   assign soundFileAmplitudes [13779] = 8'd120;
   assign soundFileAmplitudes [13780] = 8'd132;
   assign soundFileAmplitudes [13781] = 8'd144;
   assign soundFileAmplitudes [13782] = 8'd155;
   assign soundFileAmplitudes [13783] = 8'd162;
   assign soundFileAmplitudes [13784] = 8'd144;
   assign soundFileAmplitudes [13785] = 8'd119;
   assign soundFileAmplitudes [13786] = 8'd104;
   assign soundFileAmplitudes [13787] = 8'd104;
   assign soundFileAmplitudes [13788] = 8'd112;
   assign soundFileAmplitudes [13789] = 8'd115;
   assign soundFileAmplitudes [13790] = 8'd117;
   assign soundFileAmplitudes [13791] = 8'd106;
   assign soundFileAmplitudes [13792] = 8'd99;
   assign soundFileAmplitudes [13793] = 8'd95;
   assign soundFileAmplitudes [13794] = 8'd86;
   assign soundFileAmplitudes [13795] = 8'd107;
   assign soundFileAmplitudes [13796] = 8'd125;
   assign soundFileAmplitudes [13797] = 8'd144;
   assign soundFileAmplitudes [13798] = 8'd157;
   assign soundFileAmplitudes [13799] = 8'd148;
   assign soundFileAmplitudes [13800] = 8'd146;
   assign soundFileAmplitudes [13801] = 8'd149;
   assign soundFileAmplitudes [13802] = 8'd146;
   assign soundFileAmplitudes [13803] = 8'd159;
   assign soundFileAmplitudes [13804] = 8'd158;
   assign soundFileAmplitudes [13805] = 8'd141;
   assign soundFileAmplitudes [13806] = 8'd145;
   assign soundFileAmplitudes [13807] = 8'd133;
   assign soundFileAmplitudes [13808] = 8'd135;
   assign soundFileAmplitudes [13809] = 8'd116;
   assign soundFileAmplitudes [13810] = 8'd96;
   assign soundFileAmplitudes [13811] = 8'd110;
   assign soundFileAmplitudes [13812] = 8'd122;
   assign soundFileAmplitudes [13813] = 8'd134;
   assign soundFileAmplitudes [13814] = 8'd128;
   assign soundFileAmplitudes [13815] = 8'd115;
   assign soundFileAmplitudes [13816] = 8'd105;
   assign soundFileAmplitudes [13817] = 8'd108;
   assign soundFileAmplitudes [13818] = 8'd121;
   assign soundFileAmplitudes [13819] = 8'd139;
   assign soundFileAmplitudes [13820] = 8'd139;
   assign soundFileAmplitudes [13821] = 8'd120;
   assign soundFileAmplitudes [13822] = 8'd102;
   assign soundFileAmplitudes [13823] = 8'd105;
   assign soundFileAmplitudes [13824] = 8'd116;
   assign soundFileAmplitudes [13825] = 8'd125;
   assign soundFileAmplitudes [13826] = 8'd124;
   assign soundFileAmplitudes [13827] = 8'd123;
   assign soundFileAmplitudes [13828] = 8'd130;
   assign soundFileAmplitudes [13829] = 8'd120;
   assign soundFileAmplitudes [13830] = 8'd108;
   assign soundFileAmplitudes [13831] = 8'd106;
   assign soundFileAmplitudes [13832] = 8'd118;
   assign soundFileAmplitudes [13833] = 8'd139;
   assign soundFileAmplitudes [13834] = 8'd138;
   assign soundFileAmplitudes [13835] = 8'd135;
   assign soundFileAmplitudes [13836] = 8'd134;
   assign soundFileAmplitudes [13837] = 8'd127;
   assign soundFileAmplitudes [13838] = 8'd129;
   assign soundFileAmplitudes [13839] = 8'd127;
   assign soundFileAmplitudes [13840] = 8'd138;
   assign soundFileAmplitudes [13841] = 8'd126;
   assign soundFileAmplitudes [13842] = 8'd130;
   assign soundFileAmplitudes [13843] = 8'd146;
   assign soundFileAmplitudes [13844] = 8'd149;
   assign soundFileAmplitudes [13845] = 8'd155;
   assign soundFileAmplitudes [13846] = 8'd126;
   assign soundFileAmplitudes [13847] = 8'd120;
   assign soundFileAmplitudes [13848] = 8'd124;
   assign soundFileAmplitudes [13849] = 8'd130;
   assign soundFileAmplitudes [13850] = 8'd130;
   assign soundFileAmplitudes [13851] = 8'd116;
   assign soundFileAmplitudes [13852] = 8'd113;
   assign soundFileAmplitudes [13853] = 8'd109;
   assign soundFileAmplitudes [13854] = 8'd115;
   assign soundFileAmplitudes [13855] = 8'd128;
   assign soundFileAmplitudes [13856] = 8'd137;
   assign soundFileAmplitudes [13857] = 8'd138;
   assign soundFileAmplitudes [13858] = 8'd137;
   assign soundFileAmplitudes [13859] = 8'd134;
   assign soundFileAmplitudes [13860] = 8'd140;
   assign soundFileAmplitudes [13861] = 8'd129;
   assign soundFileAmplitudes [13862] = 8'd114;
   assign soundFileAmplitudes [13863] = 8'd103;
   assign soundFileAmplitudes [13864] = 8'd101;
   assign soundFileAmplitudes [13865] = 8'd115;
   assign soundFileAmplitudes [13866] = 8'd116;
   assign soundFileAmplitudes [13867] = 8'd114;
   assign soundFileAmplitudes [13868] = 8'd107;
   assign soundFileAmplitudes [13869] = 8'd104;
   assign soundFileAmplitudes [13870] = 8'd114;
   assign soundFileAmplitudes [13871] = 8'd123;
   assign soundFileAmplitudes [13872] = 8'd136;
   assign soundFileAmplitudes [13873] = 8'd134;
   assign soundFileAmplitudes [13874] = 8'd130;
   assign soundFileAmplitudes [13875] = 8'd141;
   assign soundFileAmplitudes [13876] = 8'd132;
   assign soundFileAmplitudes [13877] = 8'd127;
   assign soundFileAmplitudes [13878] = 8'd132;
   assign soundFileAmplitudes [13879] = 8'd134;
   assign soundFileAmplitudes [13880] = 8'd142;
   assign soundFileAmplitudes [13881] = 8'd146;
   assign soundFileAmplitudes [13882] = 8'd135;
   assign soundFileAmplitudes [13883] = 8'd118;
   assign soundFileAmplitudes [13884] = 8'd103;
   assign soundFileAmplitudes [13885] = 8'd93;
   assign soundFileAmplitudes [13886] = 8'd110;
   assign soundFileAmplitudes [13887] = 8'd132;
   assign soundFileAmplitudes [13888] = 8'd132;
   assign soundFileAmplitudes [13889] = 8'd128;
   assign soundFileAmplitudes [13890] = 8'd113;
   assign soundFileAmplitudes [13891] = 8'd111;
   assign soundFileAmplitudes [13892] = 8'd122;
   assign soundFileAmplitudes [13893] = 8'd141;
   assign soundFileAmplitudes [13894] = 8'd156;
   assign soundFileAmplitudes [13895] = 8'd153;
   assign soundFileAmplitudes [13896] = 8'd139;
   assign soundFileAmplitudes [13897] = 8'd116;
   assign soundFileAmplitudes [13898] = 8'd116;
   assign soundFileAmplitudes [13899] = 8'd122;
   assign soundFileAmplitudes [13900] = 8'd133;
   assign soundFileAmplitudes [13901] = 8'd141;
   assign soundFileAmplitudes [13902] = 8'd150;
   assign soundFileAmplitudes [13903] = 8'd133;
   assign soundFileAmplitudes [13904] = 8'd113;
   assign soundFileAmplitudes [13905] = 8'd107;
   assign soundFileAmplitudes [13906] = 8'd104;
   assign soundFileAmplitudes [13907] = 8'd119;
   assign soundFileAmplitudes [13908] = 8'd131;
   assign soundFileAmplitudes [13909] = 8'd140;
   assign soundFileAmplitudes [13910] = 8'd129;
   assign soundFileAmplitudes [13911] = 8'd115;
   assign soundFileAmplitudes [13912] = 8'd115;
   assign soundFileAmplitudes [13913] = 8'd111;
   assign soundFileAmplitudes [13914] = 8'd130;
   assign soundFileAmplitudes [13915] = 8'd146;
   assign soundFileAmplitudes [13916] = 8'd135;
   assign soundFileAmplitudes [13917] = 8'd137;
   assign soundFileAmplitudes [13918] = 8'd130;
   assign soundFileAmplitudes [13919] = 8'd128;
   assign soundFileAmplitudes [13920] = 8'd126;
   assign soundFileAmplitudes [13921] = 8'd115;
   assign soundFileAmplitudes [13922] = 8'd111;
   assign soundFileAmplitudes [13923] = 8'd117;
   assign soundFileAmplitudes [13924] = 8'd114;
   assign soundFileAmplitudes [13925] = 8'd102;
   assign soundFileAmplitudes [13926] = 8'd103;
   assign soundFileAmplitudes [13927] = 8'd101;
   assign soundFileAmplitudes [13928] = 8'd106;
   assign soundFileAmplitudes [13929] = 8'd122;
   assign soundFileAmplitudes [13930] = 8'd134;
   assign soundFileAmplitudes [13931] = 8'd141;
   assign soundFileAmplitudes [13932] = 8'd145;
   assign soundFileAmplitudes [13933] = 8'd130;
   assign soundFileAmplitudes [13934] = 8'd116;
   assign soundFileAmplitudes [13935] = 8'd122;
   assign soundFileAmplitudes [13936] = 8'd141;
   assign soundFileAmplitudes [13937] = 8'd158;
   assign soundFileAmplitudes [13938] = 8'd158;
   assign soundFileAmplitudes [13939] = 8'd140;
   assign soundFileAmplitudes [13940] = 8'd125;
   assign soundFileAmplitudes [13941] = 8'd123;
   assign soundFileAmplitudes [13942] = 8'd121;
   assign soundFileAmplitudes [13943] = 8'd129;
   assign soundFileAmplitudes [13944] = 8'd127;
   assign soundFileAmplitudes [13945] = 8'd130;
   assign soundFileAmplitudes [13946] = 8'd136;
   assign soundFileAmplitudes [13947] = 8'd126;
   assign soundFileAmplitudes [13948] = 8'd124;
   assign soundFileAmplitudes [13949] = 8'd127;
   assign soundFileAmplitudes [13950] = 8'd118;
   assign soundFileAmplitudes [13951] = 8'd111;
   assign soundFileAmplitudes [13952] = 8'd118;
   assign soundFileAmplitudes [13953] = 8'd117;
   assign soundFileAmplitudes [13954] = 8'd112;
   assign soundFileAmplitudes [13955] = 8'd106;
   assign soundFileAmplitudes [13956] = 8'd106;
   assign soundFileAmplitudes [13957] = 8'd128;
   assign soundFileAmplitudes [13958] = 8'd139;
   assign soundFileAmplitudes [13959] = 8'd130;
   assign soundFileAmplitudes [13960] = 8'd110;
   assign soundFileAmplitudes [13961] = 8'd101;
   assign soundFileAmplitudes [13962] = 8'd116;
   assign soundFileAmplitudes [13963] = 8'd125;
   assign soundFileAmplitudes [13964] = 8'd131;
   assign soundFileAmplitudes [13965] = 8'd127;
   assign soundFileAmplitudes [13966] = 8'd123;
   assign soundFileAmplitudes [13967] = 8'd133;
   assign soundFileAmplitudes [13968] = 8'd145;
   assign soundFileAmplitudes [13969] = 8'd144;
   assign soundFileAmplitudes [13970] = 8'd143;
   assign soundFileAmplitudes [13971] = 8'd147;
   assign soundFileAmplitudes [13972] = 8'd147;
   assign soundFileAmplitudes [13973] = 8'd151;
   assign soundFileAmplitudes [13974] = 8'd148;
   assign soundFileAmplitudes [13975] = 8'd155;
   assign soundFileAmplitudes [13976] = 8'd142;
   assign soundFileAmplitudes [13977] = 8'd132;
   assign soundFileAmplitudes [13978] = 8'd134;
   assign soundFileAmplitudes [13979] = 8'd115;
   assign soundFileAmplitudes [13980] = 8'd107;
   assign soundFileAmplitudes [13981] = 8'd107;
   assign soundFileAmplitudes [13982] = 8'd120;
   assign soundFileAmplitudes [13983] = 8'd128;
   assign soundFileAmplitudes [13984] = 8'd118;
   assign soundFileAmplitudes [13985] = 8'd119;
   assign soundFileAmplitudes [13986] = 8'd115;
   assign soundFileAmplitudes [13987] = 8'd108;
   assign soundFileAmplitudes [13988] = 8'd106;
   assign soundFileAmplitudes [13989] = 8'd113;
   assign soundFileAmplitudes [13990] = 8'd126;
   assign soundFileAmplitudes [13991] = 8'd124;
   assign soundFileAmplitudes [13992] = 8'd126;
   assign soundFileAmplitudes [13993] = 8'd116;
   assign soundFileAmplitudes [13994] = 8'd107;
   assign soundFileAmplitudes [13995] = 8'd102;
   assign soundFileAmplitudes [13996] = 8'd101;
   assign soundFileAmplitudes [13997] = 8'd91;
   assign soundFileAmplitudes [13998] = 8'd79;
   assign soundFileAmplitudes [13999] = 8'd95;
   assign soundFileAmplitudes [14000] = 8'd110;
   assign soundFileAmplitudes [14001] = 8'd119;
   assign soundFileAmplitudes [14002] = 8'd116;
   assign soundFileAmplitudes [14003] = 8'd119;
   assign soundFileAmplitudes [14004] = 8'd133;
   assign soundFileAmplitudes [14005] = 8'd152;
   assign soundFileAmplitudes [14006] = 8'd159;
   assign soundFileAmplitudes [14007] = 8'd157;
   assign soundFileAmplitudes [14008] = 8'd155;
   assign soundFileAmplitudes [14009] = 8'd151;
   assign soundFileAmplitudes [14010] = 8'd153;
   assign soundFileAmplitudes [14011] = 8'd163;
   assign soundFileAmplitudes [14012] = 8'd164;
   assign soundFileAmplitudes [14013] = 8'd155;
   assign soundFileAmplitudes [14014] = 8'd149;
   assign soundFileAmplitudes [14015] = 8'd127;
   assign soundFileAmplitudes [14016] = 8'd114;
   assign soundFileAmplitudes [14017] = 8'd122;
   assign soundFileAmplitudes [14018] = 8'd134;
   assign soundFileAmplitudes [14019] = 8'd144;
   assign soundFileAmplitudes [14020] = 8'd134;
   assign soundFileAmplitudes [14021] = 8'd124;
   assign soundFileAmplitudes [14022] = 8'd115;
   assign soundFileAmplitudes [14023] = 8'd110;
   assign soundFileAmplitudes [14024] = 8'd111;
   assign soundFileAmplitudes [14025] = 8'd116;
   assign soundFileAmplitudes [14026] = 8'd129;
   assign soundFileAmplitudes [14027] = 8'd129;
   assign soundFileAmplitudes [14028] = 8'd122;
   assign soundFileAmplitudes [14029] = 8'd109;
   assign soundFileAmplitudes [14030] = 8'd106;
   assign soundFileAmplitudes [14031] = 8'd111;
   assign soundFileAmplitudes [14032] = 8'd113;
   assign soundFileAmplitudes [14033] = 8'd111;
   assign soundFileAmplitudes [14034] = 8'd112;
   assign soundFileAmplitudes [14035] = 8'd109;
   assign soundFileAmplitudes [14036] = 8'd104;
   assign soundFileAmplitudes [14037] = 8'd109;
   assign soundFileAmplitudes [14038] = 8'd104;
   assign soundFileAmplitudes [14039] = 8'd106;
   assign soundFileAmplitudes [14040] = 8'd122;
   assign soundFileAmplitudes [14041] = 8'd134;
   assign soundFileAmplitudes [14042] = 8'd142;
   assign soundFileAmplitudes [14043] = 8'd142;
   assign soundFileAmplitudes [14044] = 8'd135;
   assign soundFileAmplitudes [14045] = 8'd146;
   assign soundFileAmplitudes [14046] = 8'd155;
   assign soundFileAmplitudes [14047] = 8'd152;
   assign soundFileAmplitudes [14048] = 8'd148;
   assign soundFileAmplitudes [14049] = 8'd137;
   assign soundFileAmplitudes [14050] = 8'd141;
   assign soundFileAmplitudes [14051] = 8'd129;
   assign soundFileAmplitudes [14052] = 8'd121;
   assign soundFileAmplitudes [14053] = 8'd122;
   assign soundFileAmplitudes [14054] = 8'd121;
   assign soundFileAmplitudes [14055] = 8'd138;
   assign soundFileAmplitudes [14056] = 8'd139;
   assign soundFileAmplitudes [14057] = 8'd125;
   assign soundFileAmplitudes [14058] = 8'd119;
   assign soundFileAmplitudes [14059] = 8'd115;
   assign soundFileAmplitudes [14060] = 8'd123;
   assign soundFileAmplitudes [14061] = 8'd142;
   assign soundFileAmplitudes [14062] = 8'd145;
   assign soundFileAmplitudes [14063] = 8'd136;
   assign soundFileAmplitudes [14064] = 8'd111;
   assign soundFileAmplitudes [14065] = 8'd95;
   assign soundFileAmplitudes [14066] = 8'd97;
   assign soundFileAmplitudes [14067] = 8'd100;
   assign soundFileAmplitudes [14068] = 8'd117;
   assign soundFileAmplitudes [14069] = 8'd127;
   assign soundFileAmplitudes [14070] = 8'd126;
   assign soundFileAmplitudes [14071] = 8'd112;
   assign soundFileAmplitudes [14072] = 8'd107;
   assign soundFileAmplitudes [14073] = 8'd111;
   assign soundFileAmplitudes [14074] = 8'd122;
   assign soundFileAmplitudes [14075] = 8'd138;
   assign soundFileAmplitudes [14076] = 8'd145;
   assign soundFileAmplitudes [14077] = 8'd151;
   assign soundFileAmplitudes [14078] = 8'd146;
   assign soundFileAmplitudes [14079] = 8'd133;
   assign soundFileAmplitudes [14080] = 8'd126;
   assign soundFileAmplitudes [14081] = 8'd124;
   assign soundFileAmplitudes [14082] = 8'd131;
   assign soundFileAmplitudes [14083] = 8'd131;
   assign soundFileAmplitudes [14084] = 8'd128;
   assign soundFileAmplitudes [14085] = 8'd127;
   assign soundFileAmplitudes [14086] = 8'd113;
   assign soundFileAmplitudes [14087] = 8'd110;
   assign soundFileAmplitudes [14088] = 8'd110;
   assign soundFileAmplitudes [14089] = 8'd120;
   assign soundFileAmplitudes [14090] = 8'd135;
   assign soundFileAmplitudes [14091] = 8'd142;
   assign soundFileAmplitudes [14092] = 8'd142;
   assign soundFileAmplitudes [14093] = 8'd134;
   assign soundFileAmplitudes [14094] = 8'd133;
   assign soundFileAmplitudes [14095] = 8'd132;
   assign soundFileAmplitudes [14096] = 8'd147;
   assign soundFileAmplitudes [14097] = 8'd146;
   assign soundFileAmplitudes [14098] = 8'd132;
   assign soundFileAmplitudes [14099] = 8'd122;
   assign soundFileAmplitudes [14100] = 8'd109;
   assign soundFileAmplitudes [14101] = 8'd100;
   assign soundFileAmplitudes [14102] = 8'd92;
   assign soundFileAmplitudes [14103] = 8'd92;
   assign soundFileAmplitudes [14104] = 8'd94;
   assign soundFileAmplitudes [14105] = 8'd104;
   assign soundFileAmplitudes [14106] = 8'd103;
   assign soundFileAmplitudes [14107] = 8'd95;
   assign soundFileAmplitudes [14108] = 8'd98;
   assign soundFileAmplitudes [14109] = 8'd115;
   assign soundFileAmplitudes [14110] = 8'd138;
   assign soundFileAmplitudes [14111] = 8'd151;
   assign soundFileAmplitudes [14112] = 8'd153;
   assign soundFileAmplitudes [14113] = 8'd155;
   assign soundFileAmplitudes [14114] = 8'd147;
   assign soundFileAmplitudes [14115] = 8'd140;
   assign soundFileAmplitudes [14116] = 8'd135;
   assign soundFileAmplitudes [14117] = 8'd133;
   assign soundFileAmplitudes [14118] = 8'd146;
   assign soundFileAmplitudes [14119] = 8'd147;
   assign soundFileAmplitudes [14120] = 8'd131;
   assign soundFileAmplitudes [14121] = 8'd118;
   assign soundFileAmplitudes [14122] = 8'd110;
   assign soundFileAmplitudes [14123] = 8'd109;
   assign soundFileAmplitudes [14124] = 8'd125;
   assign soundFileAmplitudes [14125] = 8'd148;
   assign soundFileAmplitudes [14126] = 8'd155;
   assign soundFileAmplitudes [14127] = 8'd146;
   assign soundFileAmplitudes [14128] = 8'd127;
   assign soundFileAmplitudes [14129] = 8'd120;
   assign soundFileAmplitudes [14130] = 8'd135;
   assign soundFileAmplitudes [14131] = 8'd141;
   assign soundFileAmplitudes [14132] = 8'd149;
   assign soundFileAmplitudes [14133] = 8'd140;
   assign soundFileAmplitudes [14134] = 8'd132;
   assign soundFileAmplitudes [14135] = 8'd125;
   assign soundFileAmplitudes [14136] = 8'd109;
   assign soundFileAmplitudes [14137] = 8'd96;
   assign soundFileAmplitudes [14138] = 8'd94;
   assign soundFileAmplitudes [14139] = 8'd100;
   assign soundFileAmplitudes [14140] = 8'd108;
   assign soundFileAmplitudes [14141] = 8'd117;
   assign soundFileAmplitudes [14142] = 8'd106;
   assign soundFileAmplitudes [14143] = 8'd102;
   assign soundFileAmplitudes [14144] = 8'd103;
   assign soundFileAmplitudes [14145] = 8'd125;
   assign soundFileAmplitudes [14146] = 8'd141;
   assign soundFileAmplitudes [14147] = 8'd145;
   assign soundFileAmplitudes [14148] = 8'd144;
   assign soundFileAmplitudes [14149] = 8'd141;
   assign soundFileAmplitudes [14150] = 8'd146;
   assign soundFileAmplitudes [14151] = 8'd134;
   assign soundFileAmplitudes [14152] = 8'd134;
   assign soundFileAmplitudes [14153] = 8'd136;
   assign soundFileAmplitudes [14154] = 8'd129;
   assign soundFileAmplitudes [14155] = 8'd126;
   assign soundFileAmplitudes [14156] = 8'd120;
   assign soundFileAmplitudes [14157] = 8'd112;
   assign soundFileAmplitudes [14158] = 8'd99;
   assign soundFileAmplitudes [14159] = 8'd98;
   assign soundFileAmplitudes [14160] = 8'd128;
   assign soundFileAmplitudes [14161] = 8'd149;
   assign soundFileAmplitudes [14162] = 8'd141;
   assign soundFileAmplitudes [14163] = 8'd125;
   assign soundFileAmplitudes [14164] = 8'd111;
   assign soundFileAmplitudes [14165] = 8'd126;
   assign soundFileAmplitudes [14166] = 8'd150;
   assign soundFileAmplitudes [14167] = 8'd135;
   assign soundFileAmplitudes [14168] = 8'd128;
   assign soundFileAmplitudes [14169] = 8'd121;
   assign soundFileAmplitudes [14170] = 8'd100;
   assign soundFileAmplitudes [14171] = 8'd109;
   assign soundFileAmplitudes [14172] = 8'd106;
   assign soundFileAmplitudes [14173] = 8'd114;
   assign soundFileAmplitudes [14174] = 8'd113;
   assign soundFileAmplitudes [14175] = 8'd99;
   assign soundFileAmplitudes [14176] = 8'd99;
   assign soundFileAmplitudes [14177] = 8'd100;
   assign soundFileAmplitudes [14178] = 8'd111;
   assign soundFileAmplitudes [14179] = 8'd128;
   assign soundFileAmplitudes [14180] = 8'd151;
   assign soundFileAmplitudes [14181] = 8'd163;
   assign soundFileAmplitudes [14182] = 8'd171;
   assign soundFileAmplitudes [14183] = 8'd168;
   assign soundFileAmplitudes [14184] = 8'd168;
   assign soundFileAmplitudes [14185] = 8'd172;
   assign soundFileAmplitudes [14186] = 8'd159;
   assign soundFileAmplitudes [14187] = 8'd152;
   assign soundFileAmplitudes [14188] = 8'd145;
   assign soundFileAmplitudes [14189] = 8'd130;
   assign soundFileAmplitudes [14190] = 8'd119;
   assign soundFileAmplitudes [14191] = 8'd116;
   assign soundFileAmplitudes [14192] = 8'd103;
   assign soundFileAmplitudes [14193] = 8'd96;
   assign soundFileAmplitudes [14194] = 8'd94;
   assign soundFileAmplitudes [14195] = 8'd100;
   assign soundFileAmplitudes [14196] = 8'd109;
   assign soundFileAmplitudes [14197] = 8'd111;
   assign soundFileAmplitudes [14198] = 8'd112;
   assign soundFileAmplitudes [14199] = 8'd113;
   assign soundFileAmplitudes [14200] = 8'd137;
   assign soundFileAmplitudes [14201] = 8'd152;
   assign soundFileAmplitudes [14202] = 8'd146;
   assign soundFileAmplitudes [14203] = 8'd132;
   assign soundFileAmplitudes [14204] = 8'd112;
   assign soundFileAmplitudes [14205] = 8'd93;
   assign soundFileAmplitudes [14206] = 8'd89;
   assign soundFileAmplitudes [14207] = 8'd92;
   assign soundFileAmplitudes [14208] = 8'd101;
   assign soundFileAmplitudes [14209] = 8'd112;
   assign soundFileAmplitudes [14210] = 8'd111;
   assign soundFileAmplitudes [14211] = 8'd107;
   assign soundFileAmplitudes [14212] = 8'd104;
   assign soundFileAmplitudes [14213] = 8'd118;
   assign soundFileAmplitudes [14214] = 8'd129;
   assign soundFileAmplitudes [14215] = 8'd150;
   assign soundFileAmplitudes [14216] = 8'd159;
   assign soundFileAmplitudes [14217] = 8'd169;
   assign soundFileAmplitudes [14218] = 8'd178;
   assign soundFileAmplitudes [14219] = 8'd180;
   assign soundFileAmplitudes [14220] = 8'd172;
   assign soundFileAmplitudes [14221] = 8'd158;
   assign soundFileAmplitudes [14222] = 8'd161;
   assign soundFileAmplitudes [14223] = 8'd148;
   assign soundFileAmplitudes [14224] = 8'd139;
   assign soundFileAmplitudes [14225] = 8'd123;
   assign soundFileAmplitudes [14226] = 8'd116;
   assign soundFileAmplitudes [14227] = 8'd105;
   assign soundFileAmplitudes [14228] = 8'd83;
   assign soundFileAmplitudes [14229] = 8'd80;
   assign soundFileAmplitudes [14230] = 8'd92;
   assign soundFileAmplitudes [14231] = 8'd106;
   assign soundFileAmplitudes [14232] = 8'd111;
   assign soundFileAmplitudes [14233] = 8'd108;
   assign soundFileAmplitudes [14234] = 8'd110;
   assign soundFileAmplitudes [14235] = 8'd124;
   assign soundFileAmplitudes [14236] = 8'd151;
   assign soundFileAmplitudes [14237] = 8'd144;
   assign soundFileAmplitudes [14238] = 8'd134;
   assign soundFileAmplitudes [14239] = 8'd128;
   assign soundFileAmplitudes [14240] = 8'd103;
   assign soundFileAmplitudes [14241] = 8'd113;
   assign soundFileAmplitudes [14242] = 8'd114;
   assign soundFileAmplitudes [14243] = 8'd119;
   assign soundFileAmplitudes [14244] = 8'd116;
   assign soundFileAmplitudes [14245] = 8'd111;
   assign soundFileAmplitudes [14246] = 8'd110;
   assign soundFileAmplitudes [14247] = 8'd105;
   assign soundFileAmplitudes [14248] = 8'd109;
   assign soundFileAmplitudes [14249] = 8'd116;
   assign soundFileAmplitudes [14250] = 8'd127;
   assign soundFileAmplitudes [14251] = 8'd139;
   assign soundFileAmplitudes [14252] = 8'd149;
   assign soundFileAmplitudes [14253] = 8'd151;
   assign soundFileAmplitudes [14254] = 8'd161;
   assign soundFileAmplitudes [14255] = 8'd156;
   assign soundFileAmplitudes [14256] = 8'd147;
   assign soundFileAmplitudes [14257] = 8'd146;
   assign soundFileAmplitudes [14258] = 8'd150;
   assign soundFileAmplitudes [14259] = 8'd147;
   assign soundFileAmplitudes [14260] = 8'd128;
   assign soundFileAmplitudes [14261] = 8'd114;
   assign soundFileAmplitudes [14262] = 8'd112;
   assign soundFileAmplitudes [14263] = 8'd99;
   assign soundFileAmplitudes [14264] = 8'd101;
   assign soundFileAmplitudes [14265] = 8'd124;
   assign soundFileAmplitudes [14266] = 8'd127;
   assign soundFileAmplitudes [14267] = 8'd124;
   assign soundFileAmplitudes [14268] = 8'd125;
   assign soundFileAmplitudes [14269] = 8'd124;
   assign soundFileAmplitudes [14270] = 8'd131;
   assign soundFileAmplitudes [14271] = 8'd151;
   assign soundFileAmplitudes [14272] = 8'd157;
   assign soundFileAmplitudes [14273] = 8'd143;
   assign soundFileAmplitudes [14274] = 8'd134;
   assign soundFileAmplitudes [14275] = 8'd121;
   assign soundFileAmplitudes [14276] = 8'd105;
   assign soundFileAmplitudes [14277] = 8'd95;
   assign soundFileAmplitudes [14278] = 8'd88;
   assign soundFileAmplitudes [14279] = 8'd96;
   assign soundFileAmplitudes [14280] = 8'd107;
   assign soundFileAmplitudes [14281] = 8'd100;
   assign soundFileAmplitudes [14282] = 8'd87;
   assign soundFileAmplitudes [14283] = 8'd92;
   assign soundFileAmplitudes [14284] = 8'd105;
   assign soundFileAmplitudes [14285] = 8'd126;
   assign soundFileAmplitudes [14286] = 8'd137;
   assign soundFileAmplitudes [14287] = 8'd143;
   assign soundFileAmplitudes [14288] = 8'd150;
   assign soundFileAmplitudes [14289] = 8'd159;
   assign soundFileAmplitudes [14290] = 8'd166;
   assign soundFileAmplitudes [14291] = 8'd162;
   assign soundFileAmplitudes [14292] = 8'd160;
   assign soundFileAmplitudes [14293] = 8'd160;
   assign soundFileAmplitudes [14294] = 8'd146;
   assign soundFileAmplitudes [14295] = 8'd126;
   assign soundFileAmplitudes [14296] = 8'd116;
   assign soundFileAmplitudes [14297] = 8'd105;
   assign soundFileAmplitudes [14298] = 8'd102;
   assign soundFileAmplitudes [14299] = 8'd89;
   assign soundFileAmplitudes [14300] = 8'd102;
   assign soundFileAmplitudes [14301] = 8'd113;
   assign soundFileAmplitudes [14302] = 8'd120;
   assign soundFileAmplitudes [14303] = 8'd129;
   assign soundFileAmplitudes [14304] = 8'd128;
   assign soundFileAmplitudes [14305] = 8'd132;
   assign soundFileAmplitudes [14306] = 8'd156;
   assign soundFileAmplitudes [14307] = 8'd171;
   assign soundFileAmplitudes [14308] = 8'd157;
   assign soundFileAmplitudes [14309] = 8'd152;
   assign soundFileAmplitudes [14310] = 8'd146;
   assign soundFileAmplitudes [14311] = 8'd146;
   assign soundFileAmplitudes [14312] = 8'd127;
   assign soundFileAmplitudes [14313] = 8'd116;
   assign soundFileAmplitudes [14314] = 8'd106;
   assign soundFileAmplitudes [14315] = 8'd103;
   assign soundFileAmplitudes [14316] = 8'd101;
   assign soundFileAmplitudes [14317] = 8'd91;
   assign soundFileAmplitudes [14318] = 8'd88;
   assign soundFileAmplitudes [14319] = 8'd88;
   assign soundFileAmplitudes [14320] = 8'd98;
   assign soundFileAmplitudes [14321] = 8'd113;
   assign soundFileAmplitudes [14322] = 8'd123;
   assign soundFileAmplitudes [14323] = 8'd132;
   assign soundFileAmplitudes [14324] = 8'd143;
   assign soundFileAmplitudes [14325] = 8'd153;
   assign soundFileAmplitudes [14326] = 8'd153;
   assign soundFileAmplitudes [14327] = 8'd144;
   assign soundFileAmplitudes [14328] = 8'd142;
   assign soundFileAmplitudes [14329] = 8'd135;
   assign soundFileAmplitudes [14330] = 8'd127;
   assign soundFileAmplitudes [14331] = 8'd115;
   assign soundFileAmplitudes [14332] = 8'd109;
   assign soundFileAmplitudes [14333] = 8'd95;
   assign soundFileAmplitudes [14334] = 8'd91;
   assign soundFileAmplitudes [14335] = 8'd100;
   assign soundFileAmplitudes [14336] = 8'd111;
   assign soundFileAmplitudes [14337] = 8'd120;
   assign soundFileAmplitudes [14338] = 8'd128;
   assign soundFileAmplitudes [14339] = 8'd133;
   assign soundFileAmplitudes [14340] = 8'd136;
   assign soundFileAmplitudes [14341] = 8'd145;
   assign soundFileAmplitudes [14342] = 8'd158;
   assign soundFileAmplitudes [14343] = 8'd166;
   assign soundFileAmplitudes [14344] = 8'd168;
   assign soundFileAmplitudes [14345] = 8'd172;
   assign soundFileAmplitudes [14346] = 8'd163;
   assign soundFileAmplitudes [14347] = 8'd153;
   assign soundFileAmplitudes [14348] = 8'd125;
   assign soundFileAmplitudes [14349] = 8'd114;
   assign soundFileAmplitudes [14350] = 8'd112;
   assign soundFileAmplitudes [14351] = 8'd116;
   assign soundFileAmplitudes [14352] = 8'd113;
   assign soundFileAmplitudes [14353] = 8'd99;
   assign soundFileAmplitudes [14354] = 8'd95;
   assign soundFileAmplitudes [14355] = 8'd95;
   assign soundFileAmplitudes [14356] = 8'd98;
   assign soundFileAmplitudes [14357] = 8'd102;
   assign soundFileAmplitudes [14358] = 8'd115;
   assign soundFileAmplitudes [14359] = 8'd132;
   assign soundFileAmplitudes [14360] = 8'd142;
   assign soundFileAmplitudes [14361] = 8'd136;
   assign soundFileAmplitudes [14362] = 8'd132;
   assign soundFileAmplitudes [14363] = 8'd120;
   assign soundFileAmplitudes [14364] = 8'd125;
   assign soundFileAmplitudes [14365] = 8'd125;
   assign soundFileAmplitudes [14366] = 8'd121;
   assign soundFileAmplitudes [14367] = 8'd124;
   assign soundFileAmplitudes [14368] = 8'd118;
   assign soundFileAmplitudes [14369] = 8'd108;
   assign soundFileAmplitudes [14370] = 8'd96;
   assign soundFileAmplitudes [14371] = 8'd102;
   assign soundFileAmplitudes [14372] = 8'd119;
   assign soundFileAmplitudes [14373] = 8'd135;
   assign soundFileAmplitudes [14374] = 8'd145;
   assign soundFileAmplitudes [14375] = 8'd143;
   assign soundFileAmplitudes [14376] = 8'd137;
   assign soundFileAmplitudes [14377] = 8'd131;
   assign soundFileAmplitudes [14378] = 8'd145;
   assign soundFileAmplitudes [14379] = 8'd154;
   assign soundFileAmplitudes [14380] = 8'd158;
   assign soundFileAmplitudes [14381] = 8'd157;
   assign soundFileAmplitudes [14382] = 8'd144;
   assign soundFileAmplitudes [14383] = 8'd134;
   assign soundFileAmplitudes [14384] = 8'd111;
   assign soundFileAmplitudes [14385] = 8'd103;
   assign soundFileAmplitudes [14386] = 8'd105;
   assign soundFileAmplitudes [14387] = 8'd118;
   assign soundFileAmplitudes [14388] = 8'd124;
   assign soundFileAmplitudes [14389] = 8'd126;
   assign soundFileAmplitudes [14390] = 8'd120;
   assign soundFileAmplitudes [14391] = 8'd114;
   assign soundFileAmplitudes [14392] = 8'd115;
   assign soundFileAmplitudes [14393] = 8'd116;
   assign soundFileAmplitudes [14394] = 8'd127;
   assign soundFileAmplitudes [14395] = 8'd135;
   assign soundFileAmplitudes [14396] = 8'd138;
   assign soundFileAmplitudes [14397] = 8'd135;
   assign soundFileAmplitudes [14398] = 8'd128;
   assign soundFileAmplitudes [14399] = 8'd120;
   assign soundFileAmplitudes [14400] = 8'd119;
   assign soundFileAmplitudes [14401] = 8'd112;
   assign soundFileAmplitudes [14402] = 8'd112;
   assign soundFileAmplitudes [14403] = 8'd122;
   assign soundFileAmplitudes [14404] = 8'd119;
   assign soundFileAmplitudes [14405] = 8'd96;
   assign soundFileAmplitudes [14406] = 8'd92;
   assign soundFileAmplitudes [14407] = 8'd109;
   assign soundFileAmplitudes [14408] = 8'd130;
   assign soundFileAmplitudes [14409] = 8'd145;
   assign soundFileAmplitudes [14410] = 8'd148;
   assign soundFileAmplitudes [14411] = 8'd140;
   assign soundFileAmplitudes [14412] = 8'd132;
   assign soundFileAmplitudes [14413] = 8'd138;
   assign soundFileAmplitudes [14414] = 8'd154;
   assign soundFileAmplitudes [14415] = 8'd164;
   assign soundFileAmplitudes [14416] = 8'd152;
   assign soundFileAmplitudes [14417] = 8'd151;
   assign soundFileAmplitudes [14418] = 8'd146;
   assign soundFileAmplitudes [14419] = 8'd139;
   assign soundFileAmplitudes [14420] = 8'd115;
   assign soundFileAmplitudes [14421] = 8'd95;
   assign soundFileAmplitudes [14422] = 8'd92;
   assign soundFileAmplitudes [14423] = 8'd96;
   assign soundFileAmplitudes [14424] = 8'd97;
   assign soundFileAmplitudes [14425] = 8'd103;
   assign soundFileAmplitudes [14426] = 8'd103;
   assign soundFileAmplitudes [14427] = 8'd98;
   assign soundFileAmplitudes [14428] = 8'd104;
   assign soundFileAmplitudes [14429] = 8'd113;
   assign soundFileAmplitudes [14430] = 8'd132;
   assign soundFileAmplitudes [14431] = 8'd143;
   assign soundFileAmplitudes [14432] = 8'd164;
   assign soundFileAmplitudes [14433] = 8'd161;
   assign soundFileAmplitudes [14434] = 8'd157;
   assign soundFileAmplitudes [14435] = 8'd156;
   assign soundFileAmplitudes [14436] = 8'd151;
   assign soundFileAmplitudes [14437] = 8'd155;
   assign soundFileAmplitudes [14438] = 8'd149;
   assign soundFileAmplitudes [14439] = 8'd137;
   assign soundFileAmplitudes [14440] = 8'd122;
   assign soundFileAmplitudes [14441] = 8'd105;
   assign soundFileAmplitudes [14442] = 8'd96;
   assign soundFileAmplitudes [14443] = 8'd102;
   assign soundFileAmplitudes [14444] = 8'd113;
   assign soundFileAmplitudes [14445] = 8'd126;
   assign soundFileAmplitudes [14446] = 8'd133;
   assign soundFileAmplitudes [14447] = 8'd129;
   assign soundFileAmplitudes [14448] = 8'd117;
   assign soundFileAmplitudes [14449] = 8'd107;
   assign soundFileAmplitudes [14450] = 8'd112;
   assign soundFileAmplitudes [14451] = 8'd126;
   assign soundFileAmplitudes [14452] = 8'd135;
   assign soundFileAmplitudes [14453] = 8'd136;
   assign soundFileAmplitudes [14454] = 8'd125;
   assign soundFileAmplitudes [14455] = 8'd124;
   assign soundFileAmplitudes [14456] = 8'd103;
   assign soundFileAmplitudes [14457] = 8'd81;
   assign soundFileAmplitudes [14458] = 8'd94;
   assign soundFileAmplitudes [14459] = 8'd111;
   assign soundFileAmplitudes [14460] = 8'd122;
   assign soundFileAmplitudes [14461] = 8'd124;
   assign soundFileAmplitudes [14462] = 8'd121;
   assign soundFileAmplitudes [14463] = 8'd123;
   assign soundFileAmplitudes [14464] = 8'd132;
   assign soundFileAmplitudes [14465] = 8'd139;
   assign soundFileAmplitudes [14466] = 8'd144;
   assign soundFileAmplitudes [14467] = 8'd156;
   assign soundFileAmplitudes [14468] = 8'd162;
   assign soundFileAmplitudes [14469] = 8'd155;
   assign soundFileAmplitudes [14470] = 8'd150;
   assign soundFileAmplitudes [14471] = 8'd149;
   assign soundFileAmplitudes [14472] = 8'd146;
   assign soundFileAmplitudes [14473] = 8'd143;
   assign soundFileAmplitudes [14474] = 8'd136;
   assign soundFileAmplitudes [14475] = 8'd123;
   assign soundFileAmplitudes [14476] = 8'd116;
   assign soundFileAmplitudes [14477] = 8'd102;
   assign soundFileAmplitudes [14478] = 8'd90;
   assign soundFileAmplitudes [14479] = 8'd91;
   assign soundFileAmplitudes [14480] = 8'd101;
   assign soundFileAmplitudes [14481] = 8'd118;
   assign soundFileAmplitudes [14482] = 8'd128;
   assign soundFileAmplitudes [14483] = 8'd122;
   assign soundFileAmplitudes [14484] = 8'd116;
   assign soundFileAmplitudes [14485] = 8'd117;
   assign soundFileAmplitudes [14486] = 8'd115;
   assign soundFileAmplitudes [14487] = 8'd122;
   assign soundFileAmplitudes [14488] = 8'd136;
   assign soundFileAmplitudes [14489] = 8'd148;
   assign soundFileAmplitudes [14490] = 8'd139;
   assign soundFileAmplitudes [14491] = 8'd134;
   assign soundFileAmplitudes [14492] = 8'd135;
   assign soundFileAmplitudes [14493] = 8'd125;
   assign soundFileAmplitudes [14494] = 8'd123;
   assign soundFileAmplitudes [14495] = 8'd123;
   assign soundFileAmplitudes [14496] = 8'd129;
   assign soundFileAmplitudes [14497] = 8'd131;
   assign soundFileAmplitudes [14498] = 8'd127;
   assign soundFileAmplitudes [14499] = 8'd118;
   assign soundFileAmplitudes [14500] = 8'd122;
   assign soundFileAmplitudes [14501] = 8'd125;
   assign soundFileAmplitudes [14502] = 8'd127;
   assign soundFileAmplitudes [14503] = 8'd133;
   assign soundFileAmplitudes [14504] = 8'd134;
   assign soundFileAmplitudes [14505] = 8'd138;
   assign soundFileAmplitudes [14506] = 8'd131;
   assign soundFileAmplitudes [14507] = 8'd128;
   assign soundFileAmplitudes [14508] = 8'd126;
   assign soundFileAmplitudes [14509] = 8'd124;
   assign soundFileAmplitudes [14510] = 8'd124;
   assign soundFileAmplitudes [14511] = 8'd124;
   assign soundFileAmplitudes [14512] = 8'd113;
   assign soundFileAmplitudes [14513] = 8'd102;
   assign soundFileAmplitudes [14514] = 8'd92;
   assign soundFileAmplitudes [14515] = 8'd87;
   assign soundFileAmplitudes [14516] = 8'd92;
   assign soundFileAmplitudes [14517] = 8'd105;
   assign soundFileAmplitudes [14518] = 8'd114;
   assign soundFileAmplitudes [14519] = 8'd123;
   assign soundFileAmplitudes [14520] = 8'd129;
   assign soundFileAmplitudes [14521] = 8'd137;
   assign soundFileAmplitudes [14522] = 8'd135;
   assign soundFileAmplitudes [14523] = 8'd137;
   assign soundFileAmplitudes [14524] = 8'd139;
   assign soundFileAmplitudes [14525] = 8'd144;
   assign soundFileAmplitudes [14526] = 8'd159;
   assign soundFileAmplitudes [14527] = 8'd142;
   assign soundFileAmplitudes [14528] = 8'd146;
   assign soundFileAmplitudes [14529] = 8'd140;
   assign soundFileAmplitudes [14530] = 8'd140;
   assign soundFileAmplitudes [14531] = 8'd136;
   assign soundFileAmplitudes [14532] = 8'd121;
   assign soundFileAmplitudes [14533] = 8'd129;
   assign soundFileAmplitudes [14534] = 8'd130;
   assign soundFileAmplitudes [14535] = 8'd141;
   assign soundFileAmplitudes [14536] = 8'd139;
   assign soundFileAmplitudes [14537] = 8'd131;
   assign soundFileAmplitudes [14538] = 8'd122;
   assign soundFileAmplitudes [14539] = 8'd120;
   assign soundFileAmplitudes [14540] = 8'd127;
   assign soundFileAmplitudes [14541] = 8'd127;
   assign soundFileAmplitudes [14542] = 8'd134;
   assign soundFileAmplitudes [14543] = 8'd137;
   assign soundFileAmplitudes [14544] = 8'd142;
   assign soundFileAmplitudes [14545] = 8'd138;
   assign soundFileAmplitudes [14546] = 8'd123;
   assign soundFileAmplitudes [14547] = 8'd115;
   assign soundFileAmplitudes [14548] = 8'd107;
   assign soundFileAmplitudes [14549] = 8'd104;
   assign soundFileAmplitudes [14550] = 8'd103;
   assign soundFileAmplitudes [14551] = 8'd106;
   assign soundFileAmplitudes [14552] = 8'd103;
   assign soundFileAmplitudes [14553] = 8'd91;
   assign soundFileAmplitudes [14554] = 8'd82;
   assign soundFileAmplitudes [14555] = 8'd90;
   assign soundFileAmplitudes [14556] = 8'd103;
   assign soundFileAmplitudes [14557] = 8'd117;
   assign soundFileAmplitudes [14558] = 8'd132;
   assign soundFileAmplitudes [14559] = 8'd144;
   assign soundFileAmplitudes [14560] = 8'd144;
   assign soundFileAmplitudes [14561] = 8'd135;
   assign soundFileAmplitudes [14562] = 8'd135;
   assign soundFileAmplitudes [14563] = 8'd142;
   assign soundFileAmplitudes [14564] = 8'd139;
   assign soundFileAmplitudes [14565] = 8'd151;
   assign soundFileAmplitudes [14566] = 8'd158;
   assign soundFileAmplitudes [14567] = 8'd150;
   assign soundFileAmplitudes [14568] = 8'd147;
   assign soundFileAmplitudes [14569] = 8'd118;
   assign soundFileAmplitudes [14570] = 8'd107;
   assign soundFileAmplitudes [14571] = 8'd118;
   assign soundFileAmplitudes [14572] = 8'd130;
   assign soundFileAmplitudes [14573] = 8'd130;
   assign soundFileAmplitudes [14574] = 8'd129;
   assign soundFileAmplitudes [14575] = 8'd122;
   assign soundFileAmplitudes [14576] = 8'd123;
   assign soundFileAmplitudes [14577] = 8'd122;
   assign soundFileAmplitudes [14578] = 8'd130;
   assign soundFileAmplitudes [14579] = 8'd149;
   assign soundFileAmplitudes [14580] = 8'd153;
   assign soundFileAmplitudes [14581] = 8'd158;
   assign soundFileAmplitudes [14582] = 8'd147;
   assign soundFileAmplitudes [14583] = 8'd139;
   assign soundFileAmplitudes [14584] = 8'd128;
   assign soundFileAmplitudes [14585] = 8'd124;
   assign soundFileAmplitudes [14586] = 8'd121;
   assign soundFileAmplitudes [14587] = 8'd119;
   assign soundFileAmplitudes [14588] = 8'd117;
   assign soundFileAmplitudes [14589] = 8'd113;
   assign soundFileAmplitudes [14590] = 8'd104;
   assign soundFileAmplitudes [14591] = 8'd96;
   assign soundFileAmplitudes [14592] = 8'd96;
   assign soundFileAmplitudes [14593] = 8'd103;
   assign soundFileAmplitudes [14594] = 8'd113;
   assign soundFileAmplitudes [14595] = 8'd123;
   assign soundFileAmplitudes [14596] = 8'd125;
   assign soundFileAmplitudes [14597] = 8'd118;
   assign soundFileAmplitudes [14598] = 8'd119;
   assign soundFileAmplitudes [14599] = 8'd115;
   assign soundFileAmplitudes [14600] = 8'd119;
   assign soundFileAmplitudes [14601] = 8'd136;
   assign soundFileAmplitudes [14602] = 8'd139;
   assign soundFileAmplitudes [14603] = 8'd146;
   assign soundFileAmplitudes [14604] = 8'd149;
   assign soundFileAmplitudes [14605] = 8'd141;
   assign soundFileAmplitudes [14606] = 8'd133;
   assign soundFileAmplitudes [14607] = 8'd115;
   assign soundFileAmplitudes [14608] = 8'd117;
   assign soundFileAmplitudes [14609] = 8'd117;
   assign soundFileAmplitudes [14610] = 8'd120;
   assign soundFileAmplitudes [14611] = 8'd130;
   assign soundFileAmplitudes [14612] = 8'd125;
   assign soundFileAmplitudes [14613] = 8'd120;
   assign soundFileAmplitudes [14614] = 8'd109;
   assign soundFileAmplitudes [14615] = 8'd112;
   assign soundFileAmplitudes [14616] = 8'd124;
   assign soundFileAmplitudes [14617] = 8'd137;
   assign soundFileAmplitudes [14618] = 8'd142;
   assign soundFileAmplitudes [14619] = 8'd147;
   assign soundFileAmplitudes [14620] = 8'd149;
   assign soundFileAmplitudes [14621] = 8'd147;
   assign soundFileAmplitudes [14622] = 8'd139;
   assign soundFileAmplitudes [14623] = 8'd139;
   assign soundFileAmplitudes [14624] = 8'd150;
   assign soundFileAmplitudes [14625] = 8'd144;
   assign soundFileAmplitudes [14626] = 8'd130;
   assign soundFileAmplitudes [14627] = 8'd125;
   assign soundFileAmplitudes [14628] = 8'd115;
   assign soundFileAmplitudes [14629] = 8'd92;
   assign soundFileAmplitudes [14630] = 8'd78;
   assign soundFileAmplitudes [14631] = 8'd86;
   assign soundFileAmplitudes [14632] = 8'd95;
   assign soundFileAmplitudes [14633] = 8'd108;
   assign soundFileAmplitudes [14634] = 8'd117;
   assign soundFileAmplitudes [14635] = 8'd117;
   assign soundFileAmplitudes [14636] = 8'd113;
   assign soundFileAmplitudes [14637] = 8'd112;
   assign soundFileAmplitudes [14638] = 8'd121;
   assign soundFileAmplitudes [14639] = 8'd145;
   assign soundFileAmplitudes [14640] = 8'd158;
   assign soundFileAmplitudes [14641] = 8'd154;
   assign soundFileAmplitudes [14642] = 8'd143;
   assign soundFileAmplitudes [14643] = 8'd147;
   assign soundFileAmplitudes [14644] = 8'd155;
   assign soundFileAmplitudes [14645] = 8'd125;
   assign soundFileAmplitudes [14646] = 8'd113;
   assign soundFileAmplitudes [14647] = 8'd109;
   assign soundFileAmplitudes [14648] = 8'd117;
   assign soundFileAmplitudes [14649] = 8'd126;
   assign soundFileAmplitudes [14650] = 8'd116;
   assign soundFileAmplitudes [14651] = 8'd107;
   assign soundFileAmplitudes [14652] = 8'd99;
   assign soundFileAmplitudes [14653] = 8'd102;
   assign soundFileAmplitudes [14654] = 8'd112;
   assign soundFileAmplitudes [14655] = 8'd136;
   assign soundFileAmplitudes [14656] = 8'd150;
   assign soundFileAmplitudes [14657] = 8'd163;
   assign soundFileAmplitudes [14658] = 8'd167;
   assign soundFileAmplitudes [14659] = 8'd161;
   assign soundFileAmplitudes [14660] = 8'd158;
   assign soundFileAmplitudes [14661] = 8'd152;
   assign soundFileAmplitudes [14662] = 8'd147;
   assign soundFileAmplitudes [14663] = 8'd138;
   assign soundFileAmplitudes [14664] = 8'd131;
   assign soundFileAmplitudes [14665] = 8'd119;
   assign soundFileAmplitudes [14666] = 8'd107;
   assign soundFileAmplitudes [14667] = 8'd88;
   assign soundFileAmplitudes [14668] = 8'd77;
   assign soundFileAmplitudes [14669] = 8'd83;
   assign soundFileAmplitudes [14670] = 8'd91;
   assign soundFileAmplitudes [14671] = 8'd109;
   assign soundFileAmplitudes [14672] = 8'd120;
   assign soundFileAmplitudes [14673] = 8'd127;
   assign soundFileAmplitudes [14674] = 8'd120;
   assign soundFileAmplitudes [14675] = 8'd122;
   assign soundFileAmplitudes [14676] = 8'd143;
   assign soundFileAmplitudes [14677] = 8'd145;
   assign soundFileAmplitudes [14678] = 8'd147;
   assign soundFileAmplitudes [14679] = 8'd142;
   assign soundFileAmplitudes [14680] = 8'd143;
   assign soundFileAmplitudes [14681] = 8'd142;
   assign soundFileAmplitudes [14682] = 8'd111;
   assign soundFileAmplitudes [14683] = 8'd105;
   assign soundFileAmplitudes [14684] = 8'd112;
   assign soundFileAmplitudes [14685] = 8'd120;
   assign soundFileAmplitudes [14686] = 8'd114;
   assign soundFileAmplitudes [14687] = 8'd108;
   assign soundFileAmplitudes [14688] = 8'd108;
   assign soundFileAmplitudes [14689] = 8'd112;
   assign soundFileAmplitudes [14690] = 8'd112;
   assign soundFileAmplitudes [14691] = 8'd114;
   assign soundFileAmplitudes [14692] = 8'd138;
   assign soundFileAmplitudes [14693] = 8'd151;
   assign soundFileAmplitudes [14694] = 8'd162;
   assign soundFileAmplitudes [14695] = 8'd171;
   assign soundFileAmplitudes [14696] = 8'd172;
   assign soundFileAmplitudes [14697] = 8'd165;
   assign soundFileAmplitudes [14698] = 8'd158;
   assign soundFileAmplitudes [14699] = 8'd144;
   assign soundFileAmplitudes [14700] = 8'd139;
   assign soundFileAmplitudes [14701] = 8'd123;
   assign soundFileAmplitudes [14702] = 8'd107;
   assign soundFileAmplitudes [14703] = 8'd99;
   assign soundFileAmplitudes [14704] = 8'd93;
   assign soundFileAmplitudes [14705] = 8'd96;
   assign soundFileAmplitudes [14706] = 8'd93;
   assign soundFileAmplitudes [14707] = 8'd104;
   assign soundFileAmplitudes [14708] = 8'd110;
   assign soundFileAmplitudes [14709] = 8'd116;
   assign soundFileAmplitudes [14710] = 8'd118;
   assign soundFileAmplitudes [14711] = 8'd118;
   assign soundFileAmplitudes [14712] = 8'd123;
   assign soundFileAmplitudes [14713] = 8'd139;
   assign soundFileAmplitudes [14714] = 8'd140;
   assign soundFileAmplitudes [14715] = 8'd138;
   assign soundFileAmplitudes [14716] = 8'd151;
   assign soundFileAmplitudes [14717] = 8'd149;
   assign soundFileAmplitudes [14718] = 8'd128;
   assign soundFileAmplitudes [14719] = 8'd104;
   assign soundFileAmplitudes [14720] = 8'd95;
   assign soundFileAmplitudes [14721] = 8'd104;
   assign soundFileAmplitudes [14722] = 8'd108;
   assign soundFileAmplitudes [14723] = 8'd117;
   assign soundFileAmplitudes [14724] = 8'd128;
   assign soundFileAmplitudes [14725] = 8'd123;
   assign soundFileAmplitudes [14726] = 8'd121;
   assign soundFileAmplitudes [14727] = 8'd118;
   assign soundFileAmplitudes [14728] = 8'd132;
   assign soundFileAmplitudes [14729] = 8'd152;
   assign soundFileAmplitudes [14730] = 8'd172;
   assign soundFileAmplitudes [14731] = 8'd177;
   assign soundFileAmplitudes [14732] = 8'd178;
   assign soundFileAmplitudes [14733] = 8'd170;
   assign soundFileAmplitudes [14734] = 8'd144;
   assign soundFileAmplitudes [14735] = 8'd127;
   assign soundFileAmplitudes [14736] = 8'd125;
   assign soundFileAmplitudes [14737] = 8'd124;
   assign soundFileAmplitudes [14738] = 8'd115;
   assign soundFileAmplitudes [14739] = 8'd113;
   assign soundFileAmplitudes [14740] = 8'd96;
   assign soundFileAmplitudes [14741] = 8'd85;
   assign soundFileAmplitudes [14742] = 8'd83;
   assign soundFileAmplitudes [14743] = 8'd88;
   assign soundFileAmplitudes [14744] = 8'd102;
   assign soundFileAmplitudes [14745] = 8'd118;
   assign soundFileAmplitudes [14746] = 8'd126;
   assign soundFileAmplitudes [14747] = 8'd126;
   assign soundFileAmplitudes [14748] = 8'd132;
   assign soundFileAmplitudes [14749] = 8'd135;
   assign soundFileAmplitudes [14750] = 8'd145;
   assign soundFileAmplitudes [14751] = 8'd143;
   assign soundFileAmplitudes [14752] = 8'd143;
   assign soundFileAmplitudes [14753] = 8'd139;
   assign soundFileAmplitudes [14754] = 8'd139;
   assign soundFileAmplitudes [14755] = 8'd132;
   assign soundFileAmplitudes [14756] = 8'd101;
   assign soundFileAmplitudes [14757] = 8'd95;
   assign soundFileAmplitudes [14758] = 8'd96;
   assign soundFileAmplitudes [14759] = 8'd101;
   assign soundFileAmplitudes [14760] = 8'd106;
   assign soundFileAmplitudes [14761] = 8'd102;
   assign soundFileAmplitudes [14762] = 8'd105;
   assign soundFileAmplitudes [14763] = 8'd100;
   assign soundFileAmplitudes [14764] = 8'd109;
   assign soundFileAmplitudes [14765] = 8'd132;
   assign soundFileAmplitudes [14766] = 8'd150;
   assign soundFileAmplitudes [14767] = 8'd161;
   assign soundFileAmplitudes [14768] = 8'd172;
   assign soundFileAmplitudes [14769] = 8'd171;
   assign soundFileAmplitudes [14770] = 8'd165;
   assign soundFileAmplitudes [14771] = 8'd155;
   assign soundFileAmplitudes [14772] = 8'd145;
   assign soundFileAmplitudes [14773] = 8'd137;
   assign soundFileAmplitudes [14774] = 8'd129;
   assign soundFileAmplitudes [14775] = 8'd128;
   assign soundFileAmplitudes [14776] = 8'd119;
   assign soundFileAmplitudes [14777] = 8'd114;
   assign soundFileAmplitudes [14778] = 8'd96;
   assign soundFileAmplitudes [14779] = 8'd95;
   assign soundFileAmplitudes [14780] = 8'd108;
   assign soundFileAmplitudes [14781] = 8'd122;
   assign soundFileAmplitudes [14782] = 8'd140;
   assign soundFileAmplitudes [14783] = 8'd138;
   assign soundFileAmplitudes [14784] = 8'd129;
   assign soundFileAmplitudes [14785] = 8'd118;
   assign soundFileAmplitudes [14786] = 8'd130;
   assign soundFileAmplitudes [14787] = 8'd147;
   assign soundFileAmplitudes [14788] = 8'd150;
   assign soundFileAmplitudes [14789] = 8'd149;
   assign soundFileAmplitudes [14790] = 8'd147;
   assign soundFileAmplitudes [14791] = 8'd123;
   assign soundFileAmplitudes [14792] = 8'd93;
   assign soundFileAmplitudes [14793] = 8'd72;
   assign soundFileAmplitudes [14794] = 8'd70;
   assign soundFileAmplitudes [14795] = 8'd92;
   assign soundFileAmplitudes [14796] = 8'd105;
   assign soundFileAmplitudes [14797] = 8'd105;
   assign soundFileAmplitudes [14798] = 8'd98;
   assign soundFileAmplitudes [14799] = 8'd100;
   assign soundFileAmplitudes [14800] = 8'd106;
   assign soundFileAmplitudes [14801] = 8'd122;
   assign soundFileAmplitudes [14802] = 8'd147;
   assign soundFileAmplitudes [14803] = 8'd166;
   assign soundFileAmplitudes [14804] = 8'd186;
   assign soundFileAmplitudes [14805] = 8'd191;
   assign soundFileAmplitudes [14806] = 8'd178;
   assign soundFileAmplitudes [14807] = 8'd163;
   assign soundFileAmplitudes [14808] = 8'd151;
   assign soundFileAmplitudes [14809] = 8'd149;
   assign soundFileAmplitudes [14810] = 8'd135;
   assign soundFileAmplitudes [14811] = 8'd126;
   assign soundFileAmplitudes [14812] = 8'd129;
   assign soundFileAmplitudes [14813] = 8'd123;
   assign soundFileAmplitudes [14814] = 8'd105;
   assign soundFileAmplitudes [14815] = 8'd87;
   assign soundFileAmplitudes [14816] = 8'd94;
   assign soundFileAmplitudes [14817] = 8'd109;
   assign soundFileAmplitudes [14818] = 8'd124;
   assign soundFileAmplitudes [14819] = 8'd135;
   assign soundFileAmplitudes [14820] = 8'd135;
   assign soundFileAmplitudes [14821] = 8'd126;
   assign soundFileAmplitudes [14822] = 8'd120;
   assign soundFileAmplitudes [14823] = 8'd141;
   assign soundFileAmplitudes [14824] = 8'd149;
   assign soundFileAmplitudes [14825] = 8'd131;
   assign soundFileAmplitudes [14826] = 8'd133;
   assign soundFileAmplitudes [14827] = 8'd127;
   assign soundFileAmplitudes [14828] = 8'd118;
   assign soundFileAmplitudes [14829] = 8'd96;
   assign soundFileAmplitudes [14830] = 8'd79;
   assign soundFileAmplitudes [14831] = 8'd91;
   assign soundFileAmplitudes [14832] = 8'd98;
   assign soundFileAmplitudes [14833] = 8'd94;
   assign soundFileAmplitudes [14834] = 8'd90;
   assign soundFileAmplitudes [14835] = 8'd92;
   assign soundFileAmplitudes [14836] = 8'd94;
   assign soundFileAmplitudes [14837] = 8'd104;
   assign soundFileAmplitudes [14838] = 8'd123;
   assign soundFileAmplitudes [14839] = 8'd142;
   assign soundFileAmplitudes [14840] = 8'd161;
   assign soundFileAmplitudes [14841] = 8'd178;
   assign soundFileAmplitudes [14842] = 8'd181;
   assign soundFileAmplitudes [14843] = 8'd171;
   assign soundFileAmplitudes [14844] = 8'd154;
   assign soundFileAmplitudes [14845] = 8'd149;
   assign soundFileAmplitudes [14846] = 8'd140;
   assign soundFileAmplitudes [14847] = 8'd136;
   assign soundFileAmplitudes [14848] = 8'd138;
   assign soundFileAmplitudes [14849] = 8'd128;
   assign soundFileAmplitudes [14850] = 8'd112;
   assign soundFileAmplitudes [14851] = 8'd95;
   assign soundFileAmplitudes [14852] = 8'd92;
   assign soundFileAmplitudes [14853] = 8'd105;
   assign soundFileAmplitudes [14854] = 8'd126;
   assign soundFileAmplitudes [14855] = 8'd138;
   assign soundFileAmplitudes [14856] = 8'd142;
   assign soundFileAmplitudes [14857] = 8'd124;
   assign soundFileAmplitudes [14858] = 8'd109;
   assign soundFileAmplitudes [14859] = 8'd125;
   assign soundFileAmplitudes [14860] = 8'd150;
   assign soundFileAmplitudes [14861] = 8'd154;
   assign soundFileAmplitudes [14862] = 8'd154;
   assign soundFileAmplitudes [14863] = 8'd153;
   assign soundFileAmplitudes [14864] = 8'd141;
   assign soundFileAmplitudes [14865] = 8'd128;
   assign soundFileAmplitudes [14866] = 8'd98;
   assign soundFileAmplitudes [14867] = 8'd95;
   assign soundFileAmplitudes [14868] = 8'd108;
   assign soundFileAmplitudes [14869] = 8'd116;
   assign soundFileAmplitudes [14870] = 8'd113;
   assign soundFileAmplitudes [14871] = 8'd97;
   assign soundFileAmplitudes [14872] = 8'd93;
   assign soundFileAmplitudes [14873] = 8'd95;
   assign soundFileAmplitudes [14874] = 8'd107;
   assign soundFileAmplitudes [14875] = 8'd131;
   assign soundFileAmplitudes [14876] = 8'd152;
   assign soundFileAmplitudes [14877] = 8'd166;
   assign soundFileAmplitudes [14878] = 8'd172;
   assign soundFileAmplitudes [14879] = 8'd167;
   assign soundFileAmplitudes [14880] = 8'd150;
   assign soundFileAmplitudes [14881] = 8'd138;
   assign soundFileAmplitudes [14882] = 8'd130;
   assign soundFileAmplitudes [14883] = 8'd125;
   assign soundFileAmplitudes [14884] = 8'd122;
   assign soundFileAmplitudes [14885] = 8'd115;
   assign soundFileAmplitudes [14886] = 8'd110;
   assign soundFileAmplitudes [14887] = 8'd101;
   assign soundFileAmplitudes [14888] = 8'd96;
   assign soundFileAmplitudes [14889] = 8'd98;
   assign soundFileAmplitudes [14890] = 8'd109;
   assign soundFileAmplitudes [14891] = 8'd128;
   assign soundFileAmplitudes [14892] = 8'd130;
   assign soundFileAmplitudes [14893] = 8'd132;
   assign soundFileAmplitudes [14894] = 8'd126;
   assign soundFileAmplitudes [14895] = 8'd116;
   assign soundFileAmplitudes [14896] = 8'd135;
   assign soundFileAmplitudes [14897] = 8'd149;
   assign soundFileAmplitudes [14898] = 8'd142;
   assign soundFileAmplitudes [14899] = 8'd139;
   assign soundFileAmplitudes [14900] = 8'd148;
   assign soundFileAmplitudes [14901] = 8'd148;
   assign soundFileAmplitudes [14902] = 8'd133;
   assign soundFileAmplitudes [14903] = 8'd101;
   assign soundFileAmplitudes [14904] = 8'd93;
   assign soundFileAmplitudes [14905] = 8'd102;
   assign soundFileAmplitudes [14906] = 8'd103;
   assign soundFileAmplitudes [14907] = 8'd106;
   assign soundFileAmplitudes [14908] = 8'd100;
   assign soundFileAmplitudes [14909] = 8'd97;
   assign soundFileAmplitudes [14910] = 8'd101;
   assign soundFileAmplitudes [14911] = 8'd113;
   assign soundFileAmplitudes [14912] = 8'd134;
   assign soundFileAmplitudes [14913] = 8'd157;
   assign soundFileAmplitudes [14914] = 8'd167;
   assign soundFileAmplitudes [14915] = 8'd167;
   assign soundFileAmplitudes [14916] = 8'd151;
   assign soundFileAmplitudes [14917] = 8'd148;
   assign soundFileAmplitudes [14918] = 8'd156;
   assign soundFileAmplitudes [14919] = 8'd154;
   assign soundFileAmplitudes [14920] = 8'd149;
   assign soundFileAmplitudes [14921] = 8'd131;
   assign soundFileAmplitudes [14922] = 8'd114;
   assign soundFileAmplitudes [14923] = 8'd95;
   assign soundFileAmplitudes [14924] = 8'd87;
   assign soundFileAmplitudes [14925] = 8'd84;
   assign soundFileAmplitudes [14926] = 8'd100;
   assign soundFileAmplitudes [14927] = 8'd130;
   assign soundFileAmplitudes [14928] = 8'd144;
   assign soundFileAmplitudes [14929] = 8'd139;
   assign soundFileAmplitudes [14930] = 8'd122;
   assign soundFileAmplitudes [14931] = 8'd113;
   assign soundFileAmplitudes [14932] = 8'd129;
   assign soundFileAmplitudes [14933] = 8'd153;
   assign soundFileAmplitudes [14934] = 8'd149;
   assign soundFileAmplitudes [14935] = 8'd152;
   assign soundFileAmplitudes [14936] = 8'd141;
   assign soundFileAmplitudes [14937] = 8'd136;
   assign soundFileAmplitudes [14938] = 8'd123;
   assign soundFileAmplitudes [14939] = 8'd85;
   assign soundFileAmplitudes [14940] = 8'd87;
   assign soundFileAmplitudes [14941] = 8'd97;
   assign soundFileAmplitudes [14942] = 8'd117;
   assign soundFileAmplitudes [14943] = 8'd119;
   assign soundFileAmplitudes [14944] = 8'd107;
   assign soundFileAmplitudes [14945] = 8'd107;
   assign soundFileAmplitudes [14946] = 8'd103;
   assign soundFileAmplitudes [14947] = 8'd112;
   assign soundFileAmplitudes [14948] = 8'd129;
   assign soundFileAmplitudes [14949] = 8'd148;
   assign soundFileAmplitudes [14950] = 8'd166;
   assign soundFileAmplitudes [14951] = 8'd174;
   assign soundFileAmplitudes [14952] = 8'd173;
   assign soundFileAmplitudes [14953] = 8'd161;
   assign soundFileAmplitudes [14954] = 8'd149;
   assign soundFileAmplitudes [14955] = 8'd142;
   assign soundFileAmplitudes [14956] = 8'd133;
   assign soundFileAmplitudes [14957] = 8'd120;
   assign soundFileAmplitudes [14958] = 8'd114;
   assign soundFileAmplitudes [14959] = 8'd110;
   assign soundFileAmplitudes [14960] = 8'd95;
   assign soundFileAmplitudes [14961] = 8'd87;
   assign soundFileAmplitudes [14962] = 8'd100;
   assign soundFileAmplitudes [14963] = 8'd114;
   assign soundFileAmplitudes [14964] = 8'd130;
   assign soundFileAmplitudes [14965] = 8'd134;
   assign soundFileAmplitudes [14966] = 8'd122;
   assign soundFileAmplitudes [14967] = 8'd116;
   assign soundFileAmplitudes [14968] = 8'd117;
   assign soundFileAmplitudes [14969] = 8'd124;
   assign soundFileAmplitudes [14970] = 8'd146;
   assign soundFileAmplitudes [14971] = 8'd155;
   assign soundFileAmplitudes [14972] = 8'd142;
   assign soundFileAmplitudes [14973] = 8'd140;
   assign soundFileAmplitudes [14974] = 8'd138;
   assign soundFileAmplitudes [14975] = 8'd132;
   assign soundFileAmplitudes [14976] = 8'd116;
   assign soundFileAmplitudes [14977] = 8'd99;
   assign soundFileAmplitudes [14978] = 8'd102;
   assign soundFileAmplitudes [14979] = 8'd109;
   assign soundFileAmplitudes [14980] = 8'd116;
   assign soundFileAmplitudes [14981] = 8'd113;
   assign soundFileAmplitudes [14982] = 8'd103;
   assign soundFileAmplitudes [14983] = 8'd106;
   assign soundFileAmplitudes [14984] = 8'd113;
   assign soundFileAmplitudes [14985] = 8'd139;
   assign soundFileAmplitudes [14986] = 8'd161;
   assign soundFileAmplitudes [14987] = 8'd165;
   assign soundFileAmplitudes [14988] = 8'd163;
   assign soundFileAmplitudes [14989] = 8'd152;
   assign soundFileAmplitudes [14990] = 8'd149;
   assign soundFileAmplitudes [14991] = 8'd146;
   assign soundFileAmplitudes [14992] = 8'd137;
   assign soundFileAmplitudes [14993] = 8'd129;
   assign soundFileAmplitudes [14994] = 8'd128;
   assign soundFileAmplitudes [14995] = 8'd120;
   assign soundFileAmplitudes [14996] = 8'd108;
   assign soundFileAmplitudes [14997] = 8'd98;
   assign soundFileAmplitudes [14998] = 8'd102;
   assign soundFileAmplitudes [14999] = 8'd103;
   assign soundFileAmplitudes [15000] = 8'd111;
   assign soundFileAmplitudes [15001] = 8'd113;
   assign soundFileAmplitudes [15002] = 8'd110;
   assign soundFileAmplitudes [15003] = 8'd114;
   assign soundFileAmplitudes [15004] = 8'd122;
   assign soundFileAmplitudes [15005] = 8'd127;
   assign soundFileAmplitudes [15006] = 8'd139;
   assign soundFileAmplitudes [15007] = 8'd155;
   assign soundFileAmplitudes [15008] = 8'd137;
   assign soundFileAmplitudes [15009] = 8'd137;
   assign soundFileAmplitudes [15010] = 8'd136;
   assign soundFileAmplitudes [15011] = 8'd142;
   assign soundFileAmplitudes [15012] = 8'd136;
   assign soundFileAmplitudes [15013] = 8'd105;
   assign soundFileAmplitudes [15014] = 8'd98;
   assign soundFileAmplitudes [15015] = 8'd105;
   assign soundFileAmplitudes [15016] = 8'd102;
   assign soundFileAmplitudes [15017] = 8'd104;
   assign soundFileAmplitudes [15018] = 8'd111;
   assign soundFileAmplitudes [15019] = 8'd112;
   assign soundFileAmplitudes [15020] = 8'd126;
   assign soundFileAmplitudes [15021] = 8'd141;
   assign soundFileAmplitudes [15022] = 8'd150;
   assign soundFileAmplitudes [15023] = 8'd147;
   assign soundFileAmplitudes [15024] = 8'd149;
   assign soundFileAmplitudes [15025] = 8'd148;
   assign soundFileAmplitudes [15026] = 8'd145;
   assign soundFileAmplitudes [15027] = 8'd149;
   assign soundFileAmplitudes [15028] = 8'd155;
   assign soundFileAmplitudes [15029] = 8'd152;
   assign soundFileAmplitudes [15030] = 8'd139;
   assign soundFileAmplitudes [15031] = 8'd131;
   assign soundFileAmplitudes [15032] = 8'd114;
   assign soundFileAmplitudes [15033] = 8'd107;
   assign soundFileAmplitudes [15034] = 8'd102;
   assign soundFileAmplitudes [15035] = 8'd104;
   assign soundFileAmplitudes [15036] = 8'd113;
   assign soundFileAmplitudes [15037] = 8'd123;
   assign soundFileAmplitudes [15038] = 8'd122;
   assign soundFileAmplitudes [15039] = 8'd107;
   assign soundFileAmplitudes [15040] = 8'd108;
   assign soundFileAmplitudes [15041] = 8'd111;
   assign soundFileAmplitudes [15042] = 8'd124;
   assign soundFileAmplitudes [15043] = 8'd140;
   assign soundFileAmplitudes [15044] = 8'd131;
   assign soundFileAmplitudes [15045] = 8'd133;
   assign soundFileAmplitudes [15046] = 8'd140;
   assign soundFileAmplitudes [15047] = 8'd132;
   assign soundFileAmplitudes [15048] = 8'd115;
   assign soundFileAmplitudes [15049] = 8'd87;
   assign soundFileAmplitudes [15050] = 8'd89;
   assign soundFileAmplitudes [15051] = 8'd98;
   assign soundFileAmplitudes [15052] = 8'd111;
   assign soundFileAmplitudes [15053] = 8'd126;
   assign soundFileAmplitudes [15054] = 8'd123;
   assign soundFileAmplitudes [15055] = 8'd122;
   assign soundFileAmplitudes [15056] = 8'd124;
   assign soundFileAmplitudes [15057] = 8'd138;
   assign soundFileAmplitudes [15058] = 8'd151;
   assign soundFileAmplitudes [15059] = 8'd156;
   assign soundFileAmplitudes [15060] = 8'd159;
   assign soundFileAmplitudes [15061] = 8'd159;
   assign soundFileAmplitudes [15062] = 8'd154;
   assign soundFileAmplitudes [15063] = 8'd142;
   assign soundFileAmplitudes [15064] = 8'd142;
   assign soundFileAmplitudes [15065] = 8'd149;
   assign soundFileAmplitudes [15066] = 8'd139;
   assign soundFileAmplitudes [15067] = 8'd135;
   assign soundFileAmplitudes [15068] = 8'd128;
   assign soundFileAmplitudes [15069] = 8'd111;
   assign soundFileAmplitudes [15070] = 8'd104;
   assign soundFileAmplitudes [15071] = 8'd101;
   assign soundFileAmplitudes [15072] = 8'd107;
   assign soundFileAmplitudes [15073] = 8'd124;
   assign soundFileAmplitudes [15074] = 8'd127;
   assign soundFileAmplitudes [15075] = 8'd118;
   assign soundFileAmplitudes [15076] = 8'd110;
   assign soundFileAmplitudes [15077] = 8'd113;
   assign soundFileAmplitudes [15078] = 8'd112;
   assign soundFileAmplitudes [15079] = 8'd113;
   assign soundFileAmplitudes [15080] = 8'd113;
   assign soundFileAmplitudes [15081] = 8'd112;
   assign soundFileAmplitudes [15082] = 8'd123;
   assign soundFileAmplitudes [15083] = 8'd127;
   assign soundFileAmplitudes [15084] = 8'd125;
   assign soundFileAmplitudes [15085] = 8'd102;
   assign soundFileAmplitudes [15086] = 8'd92;
   assign soundFileAmplitudes [15087] = 8'd100;
   assign soundFileAmplitudes [15088] = 8'd111;
   assign soundFileAmplitudes [15089] = 8'd123;
   assign soundFileAmplitudes [15090] = 8'd125;
   assign soundFileAmplitudes [15091] = 8'd130;
   assign soundFileAmplitudes [15092] = 8'd144;
   assign soundFileAmplitudes [15093] = 8'd155;
   assign soundFileAmplitudes [15094] = 8'd160;
   assign soundFileAmplitudes [15095] = 8'd167;
   assign soundFileAmplitudes [15096] = 8'd173;
   assign soundFileAmplitudes [15097] = 8'd163;
   assign soundFileAmplitudes [15098] = 8'd156;
   assign soundFileAmplitudes [15099] = 8'd154;
   assign soundFileAmplitudes [15100] = 8'd152;
   assign soundFileAmplitudes [15101] = 8'd143;
   assign soundFileAmplitudes [15102] = 8'd132;
   assign soundFileAmplitudes [15103] = 8'd129;
   assign soundFileAmplitudes [15104] = 8'd116;
   assign soundFileAmplitudes [15105] = 8'd103;
   assign soundFileAmplitudes [15106] = 8'd95;
   assign soundFileAmplitudes [15107] = 8'd101;
   assign soundFileAmplitudes [15108] = 8'd108;
   assign soundFileAmplitudes [15109] = 8'd123;
   assign soundFileAmplitudes [15110] = 8'd126;
   assign soundFileAmplitudes [15111] = 8'd120;
   assign soundFileAmplitudes [15112] = 8'd113;
   assign soundFileAmplitudes [15113] = 8'd112;
   assign soundFileAmplitudes [15114] = 8'd128;
   assign soundFileAmplitudes [15115] = 8'd134;
   assign soundFileAmplitudes [15116] = 8'd136;
   assign soundFileAmplitudes [15117] = 8'd129;
   assign soundFileAmplitudes [15118] = 8'd122;
   assign soundFileAmplitudes [15119] = 8'd122;
   assign soundFileAmplitudes [15120] = 8'd122;
   assign soundFileAmplitudes [15121] = 8'd112;
   assign soundFileAmplitudes [15122] = 8'd85;
   assign soundFileAmplitudes [15123] = 8'd75;
   assign soundFileAmplitudes [15124] = 8'd94;
   assign soundFileAmplitudes [15125] = 8'd114;
   assign soundFileAmplitudes [15126] = 8'd125;
   assign soundFileAmplitudes [15127] = 8'd117;
   assign soundFileAmplitudes [15128] = 8'd121;
   assign soundFileAmplitudes [15129] = 8'd136;
   assign soundFileAmplitudes [15130] = 8'd158;
   assign soundFileAmplitudes [15131] = 8'd169;
   assign soundFileAmplitudes [15132] = 8'd172;
   assign soundFileAmplitudes [15133] = 8'd167;
   assign soundFileAmplitudes [15134] = 8'd145;
   assign soundFileAmplitudes [15135] = 8'd144;
   assign soundFileAmplitudes [15136] = 8'd135;
   assign soundFileAmplitudes [15137] = 8'd131;
   assign soundFileAmplitudes [15138] = 8'd123;
   assign soundFileAmplitudes [15139] = 8'd119;
   assign soundFileAmplitudes [15140] = 8'd118;
   assign soundFileAmplitudes [15141] = 8'd110;
   assign soundFileAmplitudes [15142] = 8'd111;
   assign soundFileAmplitudes [15143] = 8'd116;
   assign soundFileAmplitudes [15144] = 8'd123;
   assign soundFileAmplitudes [15145] = 8'd133;
   assign soundFileAmplitudes [15146] = 8'd143;
   assign soundFileAmplitudes [15147] = 8'd142;
   assign soundFileAmplitudes [15148] = 8'd127;
   assign soundFileAmplitudes [15149] = 8'd118;
   assign soundFileAmplitudes [15150] = 8'd121;
   assign soundFileAmplitudes [15151] = 8'd135;
   assign soundFileAmplitudes [15152] = 8'd142;
   assign soundFileAmplitudes [15153] = 8'd134;
   assign soundFileAmplitudes [15154] = 8'd121;
   assign soundFileAmplitudes [15155] = 8'd120;
   assign soundFileAmplitudes [15156] = 8'd130;
   assign soundFileAmplitudes [15157] = 8'd119;
   assign soundFileAmplitudes [15158] = 8'd91;
   assign soundFileAmplitudes [15159] = 8'd60;
   assign soundFileAmplitudes [15160] = 8'd62;
   assign soundFileAmplitudes [15161] = 8'd84;
   assign soundFileAmplitudes [15162] = 8'd108;
   assign soundFileAmplitudes [15163] = 8'd126;
   assign soundFileAmplitudes [15164] = 8'd128;
   assign soundFileAmplitudes [15165] = 8'd140;
   assign soundFileAmplitudes [15166] = 8'd157;
   assign soundFileAmplitudes [15167] = 8'd164;
   assign soundFileAmplitudes [15168] = 8'd166;
   assign soundFileAmplitudes [15169] = 8'd159;
   assign soundFileAmplitudes [15170] = 8'd153;
   assign soundFileAmplitudes [15171] = 8'd146;
   assign soundFileAmplitudes [15172] = 8'd140;
   assign soundFileAmplitudes [15173] = 8'd139;
   assign soundFileAmplitudes [15174] = 8'd130;
   assign soundFileAmplitudes [15175] = 8'd130;
   assign soundFileAmplitudes [15176] = 8'd118;
   assign soundFileAmplitudes [15177] = 8'd119;
   assign soundFileAmplitudes [15178] = 8'd120;
   assign soundFileAmplitudes [15179] = 8'd120;
   assign soundFileAmplitudes [15180] = 8'd125;
   assign soundFileAmplitudes [15181] = 8'd127;
   assign soundFileAmplitudes [15182] = 8'd127;
   assign soundFileAmplitudes [15183] = 8'd123;
   assign soundFileAmplitudes [15184] = 8'd125;
   assign soundFileAmplitudes [15185] = 8'd118;
   assign soundFileAmplitudes [15186] = 8'd120;
   assign soundFileAmplitudes [15187] = 8'd123;
   assign soundFileAmplitudes [15188] = 8'd132;
   assign soundFileAmplitudes [15189] = 8'd126;
   assign soundFileAmplitudes [15190] = 8'd115;
   assign soundFileAmplitudes [15191] = 8'd109;
   assign soundFileAmplitudes [15192] = 8'd112;
   assign soundFileAmplitudes [15193] = 8'd107;
   assign soundFileAmplitudes [15194] = 8'd97;
   assign soundFileAmplitudes [15195] = 8'd83;
   assign soundFileAmplitudes [15196] = 8'd74;
   assign soundFileAmplitudes [15197] = 8'd93;
   assign soundFileAmplitudes [15198] = 8'd101;
   assign soundFileAmplitudes [15199] = 8'd116;
   assign soundFileAmplitudes [15200] = 8'd124;
   assign soundFileAmplitudes [15201] = 8'd133;
   assign soundFileAmplitudes [15202] = 8'd150;
   assign soundFileAmplitudes [15203] = 8'd168;
   assign soundFileAmplitudes [15204] = 8'd174;
   assign soundFileAmplitudes [15205] = 8'd174;
   assign soundFileAmplitudes [15206] = 8'd177;
   assign soundFileAmplitudes [15207] = 8'd159;
   assign soundFileAmplitudes [15208] = 8'd151;
   assign soundFileAmplitudes [15209] = 8'd145;
   assign soundFileAmplitudes [15210] = 8'd142;
   assign soundFileAmplitudes [15211] = 8'd141;
   assign soundFileAmplitudes [15212] = 8'd137;
   assign soundFileAmplitudes [15213] = 8'd134;
   assign soundFileAmplitudes [15214] = 8'd121;
   assign soundFileAmplitudes [15215] = 8'd117;
   assign soundFileAmplitudes [15216] = 8'd110;
   assign soundFileAmplitudes [15217] = 8'd108;
   assign soundFileAmplitudes [15218] = 8'd114;
   assign soundFileAmplitudes [15219] = 8'd120;
   assign soundFileAmplitudes [15220] = 8'd127;
   assign soundFileAmplitudes [15221] = 8'd126;
   assign soundFileAmplitudes [15222] = 8'd118;
   assign soundFileAmplitudes [15223] = 8'd118;
   assign soundFileAmplitudes [15224] = 8'd117;
   assign soundFileAmplitudes [15225] = 8'd111;
   assign soundFileAmplitudes [15226] = 8'd114;
   assign soundFileAmplitudes [15227] = 8'd116;
   assign soundFileAmplitudes [15228] = 8'd115;
   assign soundFileAmplitudes [15229] = 8'd117;
   assign soundFileAmplitudes [15230] = 8'd119;
   assign soundFileAmplitudes [15231] = 8'd118;
   assign soundFileAmplitudes [15232] = 8'd113;
   assign soundFileAmplitudes [15233] = 8'd97;
   assign soundFileAmplitudes [15234] = 8'd88;
   assign soundFileAmplitudes [15235] = 8'd97;
   assign soundFileAmplitudes [15236] = 8'd115;
   assign soundFileAmplitudes [15237] = 8'd134;
   assign soundFileAmplitudes [15238] = 8'd143;
   assign soundFileAmplitudes [15239] = 8'd145;
   assign soundFileAmplitudes [15240] = 8'd141;
   assign soundFileAmplitudes [15241] = 8'd141;
   assign soundFileAmplitudes [15242] = 8'd152;
   assign soundFileAmplitudes [15243] = 8'd159;
   assign soundFileAmplitudes [15244] = 8'd160;
   assign soundFileAmplitudes [15245] = 8'd158;
   assign soundFileAmplitudes [15246] = 8'd146;
   assign soundFileAmplitudes [15247] = 8'd132;
   assign soundFileAmplitudes [15248] = 8'd125;
   assign soundFileAmplitudes [15249] = 8'd129;
   assign soundFileAmplitudes [15250] = 8'd128;
   assign soundFileAmplitudes [15251] = 8'd129;
   assign soundFileAmplitudes [15252] = 8'd119;
   assign soundFileAmplitudes [15253] = 8'd108;
   assign soundFileAmplitudes [15254] = 8'd114;
   assign soundFileAmplitudes [15255] = 8'd119;
   assign soundFileAmplitudes [15256] = 8'd132;
   assign soundFileAmplitudes [15257] = 8'd133;
   assign soundFileAmplitudes [15258] = 8'd131;
   assign soundFileAmplitudes [15259] = 8'd131;
   assign soundFileAmplitudes [15260] = 8'd134;
   assign soundFileAmplitudes [15261] = 8'd135;
   assign soundFileAmplitudes [15262] = 8'd123;
   assign soundFileAmplitudes [15263] = 8'd113;
   assign soundFileAmplitudes [15264] = 8'd107;
   assign soundFileAmplitudes [15265] = 8'd107;
   assign soundFileAmplitudes [15266] = 8'd119;
   assign soundFileAmplitudes [15267] = 8'd129;
   assign soundFileAmplitudes [15268] = 8'd130;
   assign soundFileAmplitudes [15269] = 8'd118;
   assign soundFileAmplitudes [15270] = 8'd90;
   assign soundFileAmplitudes [15271] = 8'd92;
   assign soundFileAmplitudes [15272] = 8'd110;
   assign soundFileAmplitudes [15273] = 8'd124;
   assign soundFileAmplitudes [15274] = 8'd129;
   assign soundFileAmplitudes [15275] = 8'd129;
   assign soundFileAmplitudes [15276] = 8'd127;
   assign soundFileAmplitudes [15277] = 8'd137;
   assign soundFileAmplitudes [15278] = 8'd152;
   assign soundFileAmplitudes [15279] = 8'd150;
   assign soundFileAmplitudes [15280] = 8'd151;
   assign soundFileAmplitudes [15281] = 8'd143;
   assign soundFileAmplitudes [15282] = 8'd135;
   assign soundFileAmplitudes [15283] = 8'd128;
   assign soundFileAmplitudes [15284] = 8'd132;
   assign soundFileAmplitudes [15285] = 8'd130;
   assign soundFileAmplitudes [15286] = 8'd129;
   assign soundFileAmplitudes [15287] = 8'd131;
   assign soundFileAmplitudes [15288] = 8'd119;
   assign soundFileAmplitudes [15289] = 8'd111;
   assign soundFileAmplitudes [15290] = 8'd115;
   assign soundFileAmplitudes [15291] = 8'd125;
   assign soundFileAmplitudes [15292] = 8'd138;
   assign soundFileAmplitudes [15293] = 8'd144;
   assign soundFileAmplitudes [15294] = 8'd141;
   assign soundFileAmplitudes [15295] = 8'd136;
   assign soundFileAmplitudes [15296] = 8'd127;
   assign soundFileAmplitudes [15297] = 8'd121;
   assign soundFileAmplitudes [15298] = 8'd111;
   assign soundFileAmplitudes [15299] = 8'd108;
   assign soundFileAmplitudes [15300] = 8'd111;
   assign soundFileAmplitudes [15301] = 8'd109;
   assign soundFileAmplitudes [15302] = 8'd105;
   assign soundFileAmplitudes [15303] = 8'd110;
   assign soundFileAmplitudes [15304] = 8'd102;
   assign soundFileAmplitudes [15305] = 8'd102;
   assign soundFileAmplitudes [15306] = 8'd92;
   assign soundFileAmplitudes [15307] = 8'd88;
   assign soundFileAmplitudes [15308] = 8'd115;
   assign soundFileAmplitudes [15309] = 8'd133;
   assign soundFileAmplitudes [15310] = 8'd146;
   assign soundFileAmplitudes [15311] = 8'd142;
   assign soundFileAmplitudes [15312] = 8'd141;
   assign soundFileAmplitudes [15313] = 8'd137;
   assign soundFileAmplitudes [15314] = 8'd144;
   assign soundFileAmplitudes [15315] = 8'd154;
   assign soundFileAmplitudes [15316] = 8'd154;
   assign soundFileAmplitudes [15317] = 8'd151;
   assign soundFileAmplitudes [15318] = 8'd143;
   assign soundFileAmplitudes [15319] = 8'd141;
   assign soundFileAmplitudes [15320] = 8'd130;
   assign soundFileAmplitudes [15321] = 8'd130;
   assign soundFileAmplitudes [15322] = 8'd128;
   assign soundFileAmplitudes [15323] = 8'd122;
   assign soundFileAmplitudes [15324] = 8'd111;
   assign soundFileAmplitudes [15325] = 8'd98;
   assign soundFileAmplitudes [15326] = 8'd100;
   assign soundFileAmplitudes [15327] = 8'd115;
   assign soundFileAmplitudes [15328] = 8'd139;
   assign soundFileAmplitudes [15329] = 8'd147;
   assign soundFileAmplitudes [15330] = 8'd146;
   assign soundFileAmplitudes [15331] = 8'd134;
   assign soundFileAmplitudes [15332] = 8'd126;
   assign soundFileAmplitudes [15333] = 8'd129;
   assign soundFileAmplitudes [15334] = 8'd138;
   assign soundFileAmplitudes [15335] = 8'd128;
   assign soundFileAmplitudes [15336] = 8'd124;
   assign soundFileAmplitudes [15337] = 8'd122;
   assign soundFileAmplitudes [15338] = 8'd110;
   assign soundFileAmplitudes [15339] = 8'd105;
   assign soundFileAmplitudes [15340] = 8'd85;
   assign soundFileAmplitudes [15341] = 8'd83;
   assign soundFileAmplitudes [15342] = 8'd103;
   assign soundFileAmplitudes [15343] = 8'd123;
   assign soundFileAmplitudes [15344] = 8'd126;
   assign soundFileAmplitudes [15345] = 8'd123;
   assign soundFileAmplitudes [15346] = 8'd128;
   assign soundFileAmplitudes [15347] = 8'd137;
   assign soundFileAmplitudes [15348] = 8'd143;
   assign soundFileAmplitudes [15349] = 8'd154;
   assign soundFileAmplitudes [15350] = 8'd163;
   assign soundFileAmplitudes [15351] = 8'd165;
   assign soundFileAmplitudes [15352] = 8'd148;
   assign soundFileAmplitudes [15353] = 8'd133;
   assign soundFileAmplitudes [15354] = 8'd134;
   assign soundFileAmplitudes [15355] = 8'd137;
   assign soundFileAmplitudes [15356] = 8'd137;
   assign soundFileAmplitudes [15357] = 8'd133;
   assign soundFileAmplitudes [15358] = 8'd122;
   assign soundFileAmplitudes [15359] = 8'd106;
   assign soundFileAmplitudes [15360] = 8'd98;
   assign soundFileAmplitudes [15361] = 8'd97;
   assign soundFileAmplitudes [15362] = 8'd109;
   assign soundFileAmplitudes [15363] = 8'd123;
   assign soundFileAmplitudes [15364] = 8'd130;
   assign soundFileAmplitudes [15365] = 8'd128;
   assign soundFileAmplitudes [15366] = 8'd127;
   assign soundFileAmplitudes [15367] = 8'd127;
   assign soundFileAmplitudes [15368] = 8'd125;
   assign soundFileAmplitudes [15369] = 8'd126;
   assign soundFileAmplitudes [15370] = 8'd136;
   assign soundFileAmplitudes [15371] = 8'd132;
   assign soundFileAmplitudes [15372] = 8'd128;
   assign soundFileAmplitudes [15373] = 8'd123;
   assign soundFileAmplitudes [15374] = 8'd109;
   assign soundFileAmplitudes [15375] = 8'd109;
   assign soundFileAmplitudes [15376] = 8'd111;
   assign soundFileAmplitudes [15377] = 8'd123;
   assign soundFileAmplitudes [15378] = 8'd132;
   assign soundFileAmplitudes [15379] = 8'd133;
   assign soundFileAmplitudes [15380] = 8'd133;
   assign soundFileAmplitudes [15381] = 8'd130;
   assign soundFileAmplitudes [15382] = 8'd128;
   assign soundFileAmplitudes [15383] = 8'd134;
   assign soundFileAmplitudes [15384] = 8'd138;
   assign soundFileAmplitudes [15385] = 8'd140;
   assign soundFileAmplitudes [15386] = 8'd133;
   assign soundFileAmplitudes [15387] = 8'd126;
   assign soundFileAmplitudes [15388] = 8'd127;
   assign soundFileAmplitudes [15389] = 8'd125;
   assign soundFileAmplitudes [15390] = 8'd123;
   assign soundFileAmplitudes [15391] = 8'd128;
   assign soundFileAmplitudes [15392] = 8'd131;
   assign soundFileAmplitudes [15393] = 8'd119;
   assign soundFileAmplitudes [15394] = 8'd110;
   assign soundFileAmplitudes [15395] = 8'd111;
   assign soundFileAmplitudes [15396] = 8'd112;
   assign soundFileAmplitudes [15397] = 8'd119;
   assign soundFileAmplitudes [15398] = 8'd128;
   assign soundFileAmplitudes [15399] = 8'd131;
   assign soundFileAmplitudes [15400] = 8'd135;
   assign soundFileAmplitudes [15401] = 8'd139;
   assign soundFileAmplitudes [15402] = 8'd147;
   assign soundFileAmplitudes [15403] = 8'd143;
   assign soundFileAmplitudes [15404] = 8'd128;
   assign soundFileAmplitudes [15405] = 8'd117;
   assign soundFileAmplitudes [15406] = 8'd117;
   assign soundFileAmplitudes [15407] = 8'd126;
   assign soundFileAmplitudes [15408] = 8'd115;
   assign soundFileAmplitudes [15409] = 8'd116;
   assign soundFileAmplitudes [15410] = 8'd118;
   assign soundFileAmplitudes [15411] = 8'd123;
   assign soundFileAmplitudes [15412] = 8'd130;
   assign soundFileAmplitudes [15413] = 8'd122;
   assign soundFileAmplitudes [15414] = 8'd127;
   assign soundFileAmplitudes [15415] = 8'd134;
   assign soundFileAmplitudes [15416] = 8'd145;
   assign soundFileAmplitudes [15417] = 8'd147;
   assign soundFileAmplitudes [15418] = 8'd138;
   assign soundFileAmplitudes [15419] = 8'd142;
   assign soundFileAmplitudes [15420] = 8'd137;
   assign soundFileAmplitudes [15421] = 8'd135;
   assign soundFileAmplitudes [15422] = 8'd129;
   assign soundFileAmplitudes [15423] = 8'd122;
   assign soundFileAmplitudes [15424] = 8'd124;
   assign soundFileAmplitudes [15425] = 8'd124;
   assign soundFileAmplitudes [15426] = 8'd131;
   assign soundFileAmplitudes [15427] = 8'd110;
   assign soundFileAmplitudes [15428] = 8'd90;
   assign soundFileAmplitudes [15429] = 8'd90;
   assign soundFileAmplitudes [15430] = 8'd96;
   assign soundFileAmplitudes [15431] = 8'd113;
   assign soundFileAmplitudes [15432] = 8'd127;
   assign soundFileAmplitudes [15433] = 8'd135;
   assign soundFileAmplitudes [15434] = 8'd129;
   assign soundFileAmplitudes [15435] = 8'd126;
   assign soundFileAmplitudes [15436] = 8'd133;
   assign soundFileAmplitudes [15437] = 8'd133;
   assign soundFileAmplitudes [15438] = 8'd138;
   assign soundFileAmplitudes [15439] = 8'd145;
   assign soundFileAmplitudes [15440] = 8'd135;
   assign soundFileAmplitudes [15441] = 8'd133;
   assign soundFileAmplitudes [15442] = 8'd123;
   assign soundFileAmplitudes [15443] = 8'd111;
   assign soundFileAmplitudes [15444] = 8'd104;
   assign soundFileAmplitudes [15445] = 8'd95;
   assign soundFileAmplitudes [15446] = 8'd103;
   assign soundFileAmplitudes [15447] = 8'd110;
   assign soundFileAmplitudes [15448] = 8'd119;
   assign soundFileAmplitudes [15449] = 8'd130;
   assign soundFileAmplitudes [15450] = 8'd131;
   assign soundFileAmplitudes [15451] = 8'd135;
   assign soundFileAmplitudes [15452] = 8'd140;
   assign soundFileAmplitudes [15453] = 8'd145;
   assign soundFileAmplitudes [15454] = 8'd151;
   assign soundFileAmplitudes [15455] = 8'd147;
   assign soundFileAmplitudes [15456] = 8'd142;
   assign soundFileAmplitudes [15457] = 8'd133;
   assign soundFileAmplitudes [15458] = 8'd139;
   assign soundFileAmplitudes [15459] = 8'd147;
   assign soundFileAmplitudes [15460] = 8'd144;
   assign soundFileAmplitudes [15461] = 8'd140;
   assign soundFileAmplitudes [15462] = 8'd121;
   assign soundFileAmplitudes [15463] = 8'd111;
   assign soundFileAmplitudes [15464] = 8'd110;
   assign soundFileAmplitudes [15465] = 8'd112;
   assign soundFileAmplitudes [15466] = 8'd122;
   assign soundFileAmplitudes [15467] = 8'd123;
   assign soundFileAmplitudes [15468] = 8'd118;
   assign soundFileAmplitudes [15469] = 8'd109;
   assign soundFileAmplitudes [15470] = 8'd103;
   assign soundFileAmplitudes [15471] = 8'd110;
   assign soundFileAmplitudes [15472] = 8'd121;
   assign soundFileAmplitudes [15473] = 8'd127;
   assign soundFileAmplitudes [15474] = 8'd135;
   assign soundFileAmplitudes [15475] = 8'd138;
   assign soundFileAmplitudes [15476] = 8'd134;
   assign soundFileAmplitudes [15477] = 8'd130;
   assign soundFileAmplitudes [15478] = 8'd119;
   assign soundFileAmplitudes [15479] = 8'd104;
   assign soundFileAmplitudes [15480] = 8'd102;
   assign soundFileAmplitudes [15481] = 8'd121;
   assign soundFileAmplitudes [15482] = 8'd132;
   assign soundFileAmplitudes [15483] = 8'd130;
   assign soundFileAmplitudes [15484] = 8'd121;
   assign soundFileAmplitudes [15485] = 8'd110;
   assign soundFileAmplitudes [15486] = 8'd116;
   assign soundFileAmplitudes [15487] = 8'd129;
   assign soundFileAmplitudes [15488] = 8'd141;
   assign soundFileAmplitudes [15489] = 8'd149;
   assign soundFileAmplitudes [15490] = 8'd150;
   assign soundFileAmplitudes [15491] = 8'd151;
   assign soundFileAmplitudes [15492] = 8'd149;
   assign soundFileAmplitudes [15493] = 8'd147;
   assign soundFileAmplitudes [15494] = 8'd145;
   assign soundFileAmplitudes [15495] = 8'd148;
   assign soundFileAmplitudes [15496] = 8'd149;
   assign soundFileAmplitudes [15497] = 8'd135;
   assign soundFileAmplitudes [15498] = 8'd115;
   assign soundFileAmplitudes [15499] = 8'd103;
   assign soundFileAmplitudes [15500] = 8'd105;
   assign soundFileAmplitudes [15501] = 8'd117;
   assign soundFileAmplitudes [15502] = 8'd123;
   assign soundFileAmplitudes [15503] = 8'd120;
   assign soundFileAmplitudes [15504] = 8'd113;
   assign soundFileAmplitudes [15505] = 8'd109;
   assign soundFileAmplitudes [15506] = 8'd103;
   assign soundFileAmplitudes [15507] = 8'd110;
   assign soundFileAmplitudes [15508] = 8'd115;
   assign soundFileAmplitudes [15509] = 8'd108;
   assign soundFileAmplitudes [15510] = 8'd121;
   assign soundFileAmplitudes [15511] = 8'd120;
   assign soundFileAmplitudes [15512] = 8'd134;
   assign soundFileAmplitudes [15513] = 8'd129;
   assign soundFileAmplitudes [15514] = 8'd122;
   assign soundFileAmplitudes [15515] = 8'd132;
   assign soundFileAmplitudes [15516] = 8'd135;
   assign soundFileAmplitudes [15517] = 8'd137;
   assign soundFileAmplitudes [15518] = 8'd129;
   assign soundFileAmplitudes [15519] = 8'd131;
   assign soundFileAmplitudes [15520] = 8'd130;
   assign soundFileAmplitudes [15521] = 8'd140;
   assign soundFileAmplitudes [15522] = 8'd149;
   assign soundFileAmplitudes [15523] = 8'd153;
   assign soundFileAmplitudes [15524] = 8'd149;
   assign soundFileAmplitudes [15525] = 8'd137;
   assign soundFileAmplitudes [15526] = 8'd123;
   assign soundFileAmplitudes [15527] = 8'd129;
   assign soundFileAmplitudes [15528] = 8'd137;
   assign soundFileAmplitudes [15529] = 8'd138;
   assign soundFileAmplitudes [15530] = 8'd138;
   assign soundFileAmplitudes [15531] = 8'd132;
   assign soundFileAmplitudes [15532] = 8'd118;
   assign soundFileAmplitudes [15533] = 8'd98;
   assign soundFileAmplitudes [15534] = 8'd100;
   assign soundFileAmplitudes [15535] = 8'd110;
   assign soundFileAmplitudes [15536] = 8'd128;
   assign soundFileAmplitudes [15537] = 8'd142;
   assign soundFileAmplitudes [15538] = 8'd146;
   assign soundFileAmplitudes [15539] = 8'd129;
   assign soundFileAmplitudes [15540] = 8'd112;
   assign soundFileAmplitudes [15541] = 8'd114;
   assign soundFileAmplitudes [15542] = 8'd119;
   assign soundFileAmplitudes [15543] = 8'd118;
   assign soundFileAmplitudes [15544] = 8'd118;
   assign soundFileAmplitudes [15545] = 8'd121;
   assign soundFileAmplitudes [15546] = 8'd115;
   assign soundFileAmplitudes [15547] = 8'd116;
   assign soundFileAmplitudes [15548] = 8'd96;
   assign soundFileAmplitudes [15549] = 8'd100;
   assign soundFileAmplitudes [15550] = 8'd120;
   assign soundFileAmplitudes [15551] = 8'd135;
   assign soundFileAmplitudes [15552] = 8'd142;
   assign soundFileAmplitudes [15553] = 8'd134;
   assign soundFileAmplitudes [15554] = 8'd131;
   assign soundFileAmplitudes [15555] = 8'd123;
   assign soundFileAmplitudes [15556] = 8'd126;
   assign soundFileAmplitudes [15557] = 8'd130;
   assign soundFileAmplitudes [15558] = 8'd128;
   assign soundFileAmplitudes [15559] = 8'd137;
   assign soundFileAmplitudes [15560] = 8'd140;
   assign soundFileAmplitudes [15561] = 8'd136;
   assign soundFileAmplitudes [15562] = 8'd135;
   assign soundFileAmplitudes [15563] = 8'd136;
   assign soundFileAmplitudes [15564] = 8'd126;
   assign soundFileAmplitudes [15565] = 8'd119;
   assign soundFileAmplitudes [15566] = 8'd119;
   assign soundFileAmplitudes [15567] = 8'd120;
   assign soundFileAmplitudes [15568] = 8'd116;
   assign soundFileAmplitudes [15569] = 8'd113;
   assign soundFileAmplitudes [15570] = 8'd118;
   assign soundFileAmplitudes [15571] = 8'd125;
   assign soundFileAmplitudes [15572] = 8'd134;
   assign soundFileAmplitudes [15573] = 8'd137;
   assign soundFileAmplitudes [15574] = 8'd134;
   assign soundFileAmplitudes [15575] = 8'd135;
   assign soundFileAmplitudes [15576] = 8'd134;
   assign soundFileAmplitudes [15577] = 8'd136;
   assign soundFileAmplitudes [15578] = 8'd141;
   assign soundFileAmplitudes [15579] = 8'd123;
   assign soundFileAmplitudes [15580] = 8'd123;
   assign soundFileAmplitudes [15581] = 8'd126;
   assign soundFileAmplitudes [15582] = 8'd124;
   assign soundFileAmplitudes [15583] = 8'd120;
   assign soundFileAmplitudes [15584] = 8'd103;
   assign soundFileAmplitudes [15585] = 8'd103;
   assign soundFileAmplitudes [15586] = 8'd106;
   assign soundFileAmplitudes [15587] = 8'd110;
   assign soundFileAmplitudes [15588] = 8'd115;
   assign soundFileAmplitudes [15589] = 8'd125;
   assign soundFileAmplitudes [15590] = 8'd122;
   assign soundFileAmplitudes [15591] = 8'd122;
   assign soundFileAmplitudes [15592] = 8'd130;
   assign soundFileAmplitudes [15593] = 8'd136;
   assign soundFileAmplitudes [15594] = 8'd150;
   assign soundFileAmplitudes [15595] = 8'd145;
   assign soundFileAmplitudes [15596] = 8'd140;
   assign soundFileAmplitudes [15597] = 8'd143;
   assign soundFileAmplitudes [15598] = 8'd137;
   assign soundFileAmplitudes [15599] = 8'd129;
   assign soundFileAmplitudes [15600] = 8'd117;
   assign soundFileAmplitudes [15601] = 8'd114;
   assign soundFileAmplitudes [15602] = 8'd117;
   assign soundFileAmplitudes [15603] = 8'd109;
   assign soundFileAmplitudes [15604] = 8'd113;
   assign soundFileAmplitudes [15605] = 8'd118;
   assign soundFileAmplitudes [15606] = 8'd124;
   assign soundFileAmplitudes [15607] = 8'd126;
   assign soundFileAmplitudes [15608] = 8'd127;
   assign soundFileAmplitudes [15609] = 8'd126;
   assign soundFileAmplitudes [15610] = 8'd129;
   assign soundFileAmplitudes [15611] = 8'd137;
   assign soundFileAmplitudes [15612] = 8'd142;
   assign soundFileAmplitudes [15613] = 8'd151;
   assign soundFileAmplitudes [15614] = 8'd143;
   assign soundFileAmplitudes [15615] = 8'd147;
   assign soundFileAmplitudes [15616] = 8'd130;
   assign soundFileAmplitudes [15617] = 8'd130;
   assign soundFileAmplitudes [15618] = 8'd120;
   assign soundFileAmplitudes [15619] = 8'd97;
   assign soundFileAmplitudes [15620] = 8'd106;
   assign soundFileAmplitudes [15621] = 8'd109;
   assign soundFileAmplitudes [15622] = 8'd122;
   assign soundFileAmplitudes [15623] = 8'd133;
   assign soundFileAmplitudes [15624] = 8'd129;
   assign soundFileAmplitudes [15625] = 8'd127;
   assign soundFileAmplitudes [15626] = 8'd123;
   assign soundFileAmplitudes [15627] = 8'd126;
   assign soundFileAmplitudes [15628] = 8'd138;
   assign soundFileAmplitudes [15629] = 8'd144;
   assign soundFileAmplitudes [15630] = 8'd151;
   assign soundFileAmplitudes [15631] = 8'd140;
   assign soundFileAmplitudes [15632] = 8'd140;
   assign soundFileAmplitudes [15633] = 8'd136;
   assign soundFileAmplitudes [15634] = 8'd129;
   assign soundFileAmplitudes [15635] = 8'd124;
   assign soundFileAmplitudes [15636] = 8'd118;
   assign soundFileAmplitudes [15637] = 8'd115;
   assign soundFileAmplitudes [15638] = 8'd98;
   assign soundFileAmplitudes [15639] = 8'd102;
   assign soundFileAmplitudes [15640] = 8'd105;
   assign soundFileAmplitudes [15641] = 8'd107;
   assign soundFileAmplitudes [15642] = 8'd118;
   assign soundFileAmplitudes [15643] = 8'd120;
   assign soundFileAmplitudes [15644] = 8'd114;
   assign soundFileAmplitudes [15645] = 8'd108;
   assign soundFileAmplitudes [15646] = 8'd107;
   assign soundFileAmplitudes [15647] = 8'd117;
   assign soundFileAmplitudes [15648] = 8'd138;
   assign soundFileAmplitudes [15649] = 8'd137;
   assign soundFileAmplitudes [15650] = 8'd144;
   assign soundFileAmplitudes [15651] = 8'd148;
   assign soundFileAmplitudes [15652] = 8'd148;
   assign soundFileAmplitudes [15653] = 8'd145;
   assign soundFileAmplitudes [15654] = 8'd119;
   assign soundFileAmplitudes [15655] = 8'd120;
   assign soundFileAmplitudes [15656] = 8'd127;
   assign soundFileAmplitudes [15657] = 8'd142;
   assign soundFileAmplitudes [15658] = 8'd140;
   assign soundFileAmplitudes [15659] = 8'd128;
   assign soundFileAmplitudes [15660] = 8'd122;
   assign soundFileAmplitudes [15661] = 8'd116;
   assign soundFileAmplitudes [15662] = 8'd125;
   assign soundFileAmplitudes [15663] = 8'd135;
   assign soundFileAmplitudes [15664] = 8'd152;
   assign soundFileAmplitudes [15665] = 8'd160;
   assign soundFileAmplitudes [15666] = 8'd149;
   assign soundFileAmplitudes [15667] = 8'd136;
   assign soundFileAmplitudes [15668] = 8'd137;
   assign soundFileAmplitudes [15669] = 8'd139;
   assign soundFileAmplitudes [15670] = 8'd136;
   assign soundFileAmplitudes [15671] = 8'd132;
   assign soundFileAmplitudes [15672] = 8'd127;
   assign soundFileAmplitudes [15673] = 8'd116;
   assign soundFileAmplitudes [15674] = 8'd101;
   assign soundFileAmplitudes [15675] = 8'd92;
   assign soundFileAmplitudes [15676] = 8'd91;
   assign soundFileAmplitudes [15677] = 8'd101;
   assign soundFileAmplitudes [15678] = 8'd108;
   assign soundFileAmplitudes [15679] = 8'd104;
   assign soundFileAmplitudes [15680] = 8'd102;
   assign soundFileAmplitudes [15681] = 8'd109;
   assign soundFileAmplitudes [15682] = 8'd112;
   assign soundFileAmplitudes [15683] = 8'd118;
   assign soundFileAmplitudes [15684] = 8'd124;
   assign soundFileAmplitudes [15685] = 8'd127;
   assign soundFileAmplitudes [15686] = 8'd140;
   assign soundFileAmplitudes [15687] = 8'd142;
   assign soundFileAmplitudes [15688] = 8'd153;
   assign soundFileAmplitudes [15689] = 8'd140;
   assign soundFileAmplitudes [15690] = 8'd125;
   assign soundFileAmplitudes [15691] = 8'd130;
   assign soundFileAmplitudes [15692] = 8'd126;
   assign soundFileAmplitudes [15693] = 8'd132;
   assign soundFileAmplitudes [15694] = 8'd128;
   assign soundFileAmplitudes [15695] = 8'd126;
   assign soundFileAmplitudes [15696] = 8'd122;
   assign soundFileAmplitudes [15697] = 8'd128;
   assign soundFileAmplitudes [15698] = 8'd138;
   assign soundFileAmplitudes [15699] = 8'd144;
   assign soundFileAmplitudes [15700] = 8'd155;
   assign soundFileAmplitudes [15701] = 8'd152;
   assign soundFileAmplitudes [15702] = 8'd140;
   assign soundFileAmplitudes [15703] = 8'd136;
   assign soundFileAmplitudes [15704] = 8'd134;
   assign soundFileAmplitudes [15705] = 8'd130;
   assign soundFileAmplitudes [15706] = 8'd130;
   assign soundFileAmplitudes [15707] = 8'd135;
   assign soundFileAmplitudes [15708] = 8'd129;
   assign soundFileAmplitudes [15709] = 8'd106;
   assign soundFileAmplitudes [15710] = 8'd92;
   assign soundFileAmplitudes [15711] = 8'd87;
   assign soundFileAmplitudes [15712] = 8'd87;
   assign soundFileAmplitudes [15713] = 8'd100;
   assign soundFileAmplitudes [15714] = 8'd111;
   assign soundFileAmplitudes [15715] = 8'd112;
   assign soundFileAmplitudes [15716] = 8'd111;
   assign soundFileAmplitudes [15717] = 8'd109;
   assign soundFileAmplitudes [15718] = 8'd115;
   assign soundFileAmplitudes [15719] = 8'd125;
   assign soundFileAmplitudes [15720] = 8'd133;
   assign soundFileAmplitudes [15721] = 8'd142;
   assign soundFileAmplitudes [15722] = 8'd143;
   assign soundFileAmplitudes [15723] = 8'd135;
   assign soundFileAmplitudes [15724] = 8'd136;
   assign soundFileAmplitudes [15725] = 8'd119;
   assign soundFileAmplitudes [15726] = 8'd111;
   assign soundFileAmplitudes [15727] = 8'd118;
   assign soundFileAmplitudes [15728] = 8'd127;
   assign soundFileAmplitudes [15729] = 8'd134;
   assign soundFileAmplitudes [15730] = 8'd131;
   assign soundFileAmplitudes [15731] = 8'd133;
   assign soundFileAmplitudes [15732] = 8'd137;
   assign soundFileAmplitudes [15733] = 8'd149;
   assign soundFileAmplitudes [15734] = 8'd155;
   assign soundFileAmplitudes [15735] = 8'd157;
   assign soundFileAmplitudes [15736] = 8'd151;
   assign soundFileAmplitudes [15737] = 8'd140;
   assign soundFileAmplitudes [15738] = 8'd147;
   assign soundFileAmplitudes [15739] = 8'd151;
   assign soundFileAmplitudes [15740] = 8'd145;
   assign soundFileAmplitudes [15741] = 8'd135;
   assign soundFileAmplitudes [15742] = 8'd130;
   assign soundFileAmplitudes [15743] = 8'd130;
   assign soundFileAmplitudes [15744] = 8'd112;
   assign soundFileAmplitudes [15745] = 8'd95;
   assign soundFileAmplitudes [15746] = 8'd93;
   assign soundFileAmplitudes [15747] = 8'd96;
   assign soundFileAmplitudes [15748] = 8'd105;
   assign soundFileAmplitudes [15749] = 8'd108;
   assign soundFileAmplitudes [15750] = 8'd107;
   assign soundFileAmplitudes [15751] = 8'd109;
   assign soundFileAmplitudes [15752] = 8'd110;
   assign soundFileAmplitudes [15753] = 8'd116;
   assign soundFileAmplitudes [15754] = 8'd122;
   assign soundFileAmplitudes [15755] = 8'd126;
   assign soundFileAmplitudes [15756] = 8'd128;
   assign soundFileAmplitudes [15757] = 8'd126;
   assign soundFileAmplitudes [15758] = 8'd134;
   assign soundFileAmplitudes [15759] = 8'd129;
   assign soundFileAmplitudes [15760] = 8'd121;
   assign soundFileAmplitudes [15761] = 8'd113;
   assign soundFileAmplitudes [15762] = 8'd107;
   assign soundFileAmplitudes [15763] = 8'd108;
   assign soundFileAmplitudes [15764] = 8'd116;
   assign soundFileAmplitudes [15765] = 8'd132;
   assign soundFileAmplitudes [15766] = 8'd137;
   assign soundFileAmplitudes [15767] = 8'd144;
   assign soundFileAmplitudes [15768] = 8'd141;
   assign soundFileAmplitudes [15769] = 8'd143;
   assign soundFileAmplitudes [15770] = 8'd144;
   assign soundFileAmplitudes [15771] = 8'd155;
   assign soundFileAmplitudes [15772] = 8'd168;
   assign soundFileAmplitudes [15773] = 8'd159;
   assign soundFileAmplitudes [15774] = 8'd157;
   assign soundFileAmplitudes [15775] = 8'd148;
   assign soundFileAmplitudes [15776] = 8'd138;
   assign soundFileAmplitudes [15777] = 8'd135;
   assign soundFileAmplitudes [15778] = 8'd125;
   assign soundFileAmplitudes [15779] = 8'd116;
   assign soundFileAmplitudes [15780] = 8'd107;
   assign soundFileAmplitudes [15781] = 8'd104;
   assign soundFileAmplitudes [15782] = 8'd109;
   assign soundFileAmplitudes [15783] = 8'd112;
   assign soundFileAmplitudes [15784] = 8'd115;
   assign soundFileAmplitudes [15785] = 8'd109;
   assign soundFileAmplitudes [15786] = 8'd102;
   assign soundFileAmplitudes [15787] = 8'd112;
   assign soundFileAmplitudes [15788] = 8'd123;
   assign soundFileAmplitudes [15789] = 8'd128;
   assign soundFileAmplitudes [15790] = 8'd141;
   assign soundFileAmplitudes [15791] = 8'd129;
   assign soundFileAmplitudes [15792] = 8'd123;
   assign soundFileAmplitudes [15793] = 8'd126;
   assign soundFileAmplitudes [15794] = 8'd134;
   assign soundFileAmplitudes [15795] = 8'd133;
   assign soundFileAmplitudes [15796] = 8'd110;
   assign soundFileAmplitudes [15797] = 8'd117;
   assign soundFileAmplitudes [15798] = 8'd134;
   assign soundFileAmplitudes [15799] = 8'd139;
   assign soundFileAmplitudes [15800] = 8'd127;
   assign soundFileAmplitudes [15801] = 8'd112;
   assign soundFileAmplitudes [15802] = 8'd104;
   assign soundFileAmplitudes [15803] = 8'd115;
   assign soundFileAmplitudes [15804] = 8'd137;
   assign soundFileAmplitudes [15805] = 8'd153;
   assign soundFileAmplitudes [15806] = 8'd154;
   assign soundFileAmplitudes [15807] = 8'd150;
   assign soundFileAmplitudes [15808] = 8'd137;
   assign soundFileAmplitudes [15809] = 8'd136;
   assign soundFileAmplitudes [15810] = 8'd151;
   assign soundFileAmplitudes [15811] = 8'd145;
   assign soundFileAmplitudes [15812] = 8'd135;
   assign soundFileAmplitudes [15813] = 8'd124;
   assign soundFileAmplitudes [15814] = 8'd120;
   assign soundFileAmplitudes [15815] = 8'd116;
   assign soundFileAmplitudes [15816] = 8'd109;
   assign soundFileAmplitudes [15817] = 8'd103;
   assign soundFileAmplitudes [15818] = 8'd96;
   assign soundFileAmplitudes [15819] = 8'd104;
   assign soundFileAmplitudes [15820] = 8'd113;
   assign soundFileAmplitudes [15821] = 8'd120;
   assign soundFileAmplitudes [15822] = 8'd117;
   assign soundFileAmplitudes [15823] = 8'd117;
   assign soundFileAmplitudes [15824] = 8'd123;
   assign soundFileAmplitudes [15825] = 8'd131;
   assign soundFileAmplitudes [15826] = 8'd141;
   assign soundFileAmplitudes [15827] = 8'd135;
   assign soundFileAmplitudes [15828] = 8'd132;
   assign soundFileAmplitudes [15829] = 8'd129;
   assign soundFileAmplitudes [15830] = 8'd129;
   assign soundFileAmplitudes [15831] = 8'd129;
   assign soundFileAmplitudes [15832] = 8'd113;
   assign soundFileAmplitudes [15833] = 8'd109;
   assign soundFileAmplitudes [15834] = 8'd117;
   assign soundFileAmplitudes [15835] = 8'd118;
   assign soundFileAmplitudes [15836] = 8'd121;
   assign soundFileAmplitudes [15837] = 8'd125;
   assign soundFileAmplitudes [15838] = 8'd122;
   assign soundFileAmplitudes [15839] = 8'd115;
   assign soundFileAmplitudes [15840] = 8'd118;
   assign soundFileAmplitudes [15841] = 8'd130;
   assign soundFileAmplitudes [15842] = 8'd145;
   assign soundFileAmplitudes [15843] = 8'd152;
   assign soundFileAmplitudes [15844] = 8'd148;
   assign soundFileAmplitudes [15845] = 8'd138;
   assign soundFileAmplitudes [15846] = 8'd122;
   assign soundFileAmplitudes [15847] = 8'd119;
   assign soundFileAmplitudes [15848] = 8'd127;
   assign soundFileAmplitudes [15849] = 8'd137;
   assign soundFileAmplitudes [15850] = 8'd147;
   assign soundFileAmplitudes [15851] = 8'd139;
   assign soundFileAmplitudes [15852] = 8'd137;
   assign soundFileAmplitudes [15853] = 8'd140;
   assign soundFileAmplitudes [15854] = 8'd129;
   assign soundFileAmplitudes [15855] = 8'd122;
   assign soundFileAmplitudes [15856] = 8'd127;
   assign soundFileAmplitudes [15857] = 8'd134;
   assign soundFileAmplitudes [15858] = 8'd132;
   assign soundFileAmplitudes [15859] = 8'd125;
   assign soundFileAmplitudes [15860] = 8'd117;
   assign soundFileAmplitudes [15861] = 8'd114;
   assign soundFileAmplitudes [15862] = 8'd118;
   assign soundFileAmplitudes [15863] = 8'd123;
   assign soundFileAmplitudes [15864] = 8'd126;
   assign soundFileAmplitudes [15865] = 8'd129;
   assign soundFileAmplitudes [15866] = 8'd134;
   assign soundFileAmplitudes [15867] = 8'd133;
   assign soundFileAmplitudes [15868] = 8'd128;
   assign soundFileAmplitudes [15869] = 8'd124;
   assign soundFileAmplitudes [15870] = 8'd123;
   assign soundFileAmplitudes [15871] = 8'd128;
   assign soundFileAmplitudes [15872] = 8'd134;
   assign soundFileAmplitudes [15873] = 8'd128;
   assign soundFileAmplitudes [15874] = 8'd121;
   assign soundFileAmplitudes [15875] = 8'd115;
   assign soundFileAmplitudes [15876] = 8'd108;
   assign soundFileAmplitudes [15877] = 8'd114;
   assign soundFileAmplitudes [15878] = 8'd124;
   assign soundFileAmplitudes [15879] = 8'd126;
   assign soundFileAmplitudes [15880] = 8'd127;
   assign soundFileAmplitudes [15881] = 8'd124;
   assign soundFileAmplitudes [15882] = 8'd127;
   assign soundFileAmplitudes [15883] = 8'd122;
   assign soundFileAmplitudes [15884] = 8'd124;
   assign soundFileAmplitudes [15885] = 8'd139;
   assign soundFileAmplitudes [15886] = 8'd141;
   assign soundFileAmplitudes [15887] = 8'd146;
   assign soundFileAmplitudes [15888] = 8'd148;
   assign soundFileAmplitudes [15889] = 8'd154;
   assign soundFileAmplitudes [15890] = 8'd149;
   assign soundFileAmplitudes [15891] = 8'd135;
   assign soundFileAmplitudes [15892] = 8'd132;
   assign soundFileAmplitudes [15893] = 8'd129;
   assign soundFileAmplitudes [15894] = 8'd129;
   assign soundFileAmplitudes [15895] = 8'd123;
   assign soundFileAmplitudes [15896] = 8'd115;
   assign soundFileAmplitudes [15897] = 8'd117;
   assign soundFileAmplitudes [15898] = 8'd107;
   assign soundFileAmplitudes [15899] = 8'd101;
   assign soundFileAmplitudes [15900] = 8'd105;
   assign soundFileAmplitudes [15901] = 8'd112;
   assign soundFileAmplitudes [15902] = 8'd121;
   assign soundFileAmplitudes [15903] = 8'd130;
   assign soundFileAmplitudes [15904] = 8'd128;
   assign soundFileAmplitudes [15905] = 8'd124;
   assign soundFileAmplitudes [15906] = 8'd124;
   assign soundFileAmplitudes [15907] = 8'd134;
   assign soundFileAmplitudes [15908] = 8'd140;
   assign soundFileAmplitudes [15909] = 8'd132;
   assign soundFileAmplitudes [15910] = 8'd131;
   assign soundFileAmplitudes [15911] = 8'd119;
   assign soundFileAmplitudes [15912] = 8'd109;
   assign soundFileAmplitudes [15913] = 8'd101;
   assign soundFileAmplitudes [15914] = 8'd107;
   assign soundFileAmplitudes [15915] = 8'd116;
   assign soundFileAmplitudes [15916] = 8'd121;
   assign soundFileAmplitudes [15917] = 8'd125;
   assign soundFileAmplitudes [15918] = 8'd116;
   assign soundFileAmplitudes [15919] = 8'd121;
   assign soundFileAmplitudes [15920] = 8'd136;
   assign soundFileAmplitudes [15921] = 8'd148;
   assign soundFileAmplitudes [15922] = 8'd154;
   assign soundFileAmplitudes [15923] = 8'd154;
   assign soundFileAmplitudes [15924] = 8'd151;
   assign soundFileAmplitudes [15925] = 8'd148;
   assign soundFileAmplitudes [15926] = 8'd138;
   assign soundFileAmplitudes [15927] = 8'd134;
   assign soundFileAmplitudes [15928] = 8'd139;
   assign soundFileAmplitudes [15929] = 8'd134;
   assign soundFileAmplitudes [15930] = 8'd126;
   assign soundFileAmplitudes [15931] = 8'd113;
   assign soundFileAmplitudes [15932] = 8'd104;
   assign soundFileAmplitudes [15933] = 8'd101;
   assign soundFileAmplitudes [15934] = 8'd100;
   assign soundFileAmplitudes [15935] = 8'd106;
   assign soundFileAmplitudes [15936] = 8'd111;
   assign soundFileAmplitudes [15937] = 8'd113;
   assign soundFileAmplitudes [15938] = 8'd114;
   assign soundFileAmplitudes [15939] = 8'd118;
   assign soundFileAmplitudes [15940] = 8'd125;
   assign soundFileAmplitudes [15941] = 8'd134;
   assign soundFileAmplitudes [15942] = 8'd134;
   assign soundFileAmplitudes [15943] = 8'd138;
   assign soundFileAmplitudes [15944] = 8'd140;
   assign soundFileAmplitudes [15945] = 8'd136;
   assign soundFileAmplitudes [15946] = 8'd128;
   assign soundFileAmplitudes [15947] = 8'd116;
   assign soundFileAmplitudes [15948] = 8'd119;
   assign soundFileAmplitudes [15949] = 8'd115;
   assign soundFileAmplitudes [15950] = 8'd121;
   assign soundFileAmplitudes [15951] = 8'd125;
   assign soundFileAmplitudes [15952] = 8'd123;
   assign soundFileAmplitudes [15953] = 8'd124;
   assign soundFileAmplitudes [15954] = 8'd121;
   assign soundFileAmplitudes [15955] = 8'd128;
   assign soundFileAmplitudes [15956] = 8'd140;
   assign soundFileAmplitudes [15957] = 8'd146;
   assign soundFileAmplitudes [15958] = 8'd144;
   assign soundFileAmplitudes [15959] = 8'd142;
   assign soundFileAmplitudes [15960] = 8'd136;
   assign soundFileAmplitudes [15961] = 8'd132;
   assign soundFileAmplitudes [15962] = 8'd127;
   assign soundFileAmplitudes [15963] = 8'd130;
   assign soundFileAmplitudes [15964] = 8'd132;
   assign soundFileAmplitudes [15965] = 8'd125;
   assign soundFileAmplitudes [15966] = 8'd110;
   assign soundFileAmplitudes [15967] = 8'd104;
   assign soundFileAmplitudes [15968] = 8'd107;
   assign soundFileAmplitudes [15969] = 8'd112;
   assign soundFileAmplitudes [15970] = 8'd118;
   assign soundFileAmplitudes [15971] = 8'd122;
   assign soundFileAmplitudes [15972] = 8'd115;
   assign soundFileAmplitudes [15973] = 8'd121;
   assign soundFileAmplitudes [15974] = 8'd140;
   assign soundFileAmplitudes [15975] = 8'd138;
   assign soundFileAmplitudes [15976] = 8'd133;
   assign soundFileAmplitudes [15977] = 8'd133;
   assign soundFileAmplitudes [15978] = 8'd136;
   assign soundFileAmplitudes [15979] = 8'd144;
   assign soundFileAmplitudes [15980] = 8'd134;
   assign soundFileAmplitudes [15981] = 8'd110;
   assign soundFileAmplitudes [15982] = 8'd102;
   assign soundFileAmplitudes [15983] = 8'd108;
   assign soundFileAmplitudes [15984] = 8'd118;
   assign soundFileAmplitudes [15985] = 8'd128;
   assign soundFileAmplitudes [15986] = 8'd133;
   assign soundFileAmplitudes [15987] = 8'd131;
   assign soundFileAmplitudes [15988] = 8'd131;
   assign soundFileAmplitudes [15989] = 8'd127;
   assign soundFileAmplitudes [15990] = 8'd130;
   assign soundFileAmplitudes [15991] = 8'd145;
   assign soundFileAmplitudes [15992] = 8'd155;
   assign soundFileAmplitudes [15993] = 8'd156;
   assign soundFileAmplitudes [15994] = 8'd151;
   assign soundFileAmplitudes [15995] = 8'd147;
   assign soundFileAmplitudes [15996] = 8'd143;
   assign soundFileAmplitudes [15997] = 8'd127;
   assign soundFileAmplitudes [15998] = 8'd120;
   assign soundFileAmplitudes [15999] = 8'd116;
   assign soundFileAmplitudes [16000] = 8'd107;
   assign soundFileAmplitudes [16001] = 8'd113;
   assign soundFileAmplitudes [16002] = 8'd113;
   assign soundFileAmplitudes [16003] = 8'd118;
   assign soundFileAmplitudes [16004] = 8'd110;
   assign soundFileAmplitudes [16005] = 8'd94;
   assign soundFileAmplitudes [16006] = 8'd105;
   assign soundFileAmplitudes [16007] = 8'd118;
   assign soundFileAmplitudes [16008] = 8'd136;
   assign soundFileAmplitudes [16009] = 8'd147;
   assign soundFileAmplitudes [16010] = 8'd137;
   assign soundFileAmplitudes [16011] = 8'd131;
   assign soundFileAmplitudes [16012] = 8'd127;
   assign soundFileAmplitudes [16013] = 8'd125;
   assign soundFileAmplitudes [16014] = 8'd127;
   assign soundFileAmplitudes [16015] = 8'd118;
   assign soundFileAmplitudes [16016] = 8'd114;
   assign soundFileAmplitudes [16017] = 8'd115;
   assign soundFileAmplitudes [16018] = 8'd116;
   assign soundFileAmplitudes [16019] = 8'd111;
   assign soundFileAmplitudes [16020] = 8'd123;
   assign soundFileAmplitudes [16021] = 8'd139;
   assign soundFileAmplitudes [16022] = 8'd142;
   assign soundFileAmplitudes [16023] = 8'd147;
   assign soundFileAmplitudes [16024] = 8'd138;
   assign soundFileAmplitudes [16025] = 8'd135;
   assign soundFileAmplitudes [16026] = 8'd146;
   assign soundFileAmplitudes [16027] = 8'd154;
   assign soundFileAmplitudes [16028] = 8'd160;
   assign soundFileAmplitudes [16029] = 8'd154;
   assign soundFileAmplitudes [16030] = 8'd142;
   assign soundFileAmplitudes [16031] = 8'd132;
   assign soundFileAmplitudes [16032] = 8'd113;
   assign soundFileAmplitudes [16033] = 8'd107;
   assign soundFileAmplitudes [16034] = 8'd108;
   assign soundFileAmplitudes [16035] = 8'd110;
   assign soundFileAmplitudes [16036] = 8'd111;
   assign soundFileAmplitudes [16037] = 8'd106;
   assign soundFileAmplitudes [16038] = 8'd108;
   assign soundFileAmplitudes [16039] = 8'd116;
   assign soundFileAmplitudes [16040] = 8'd118;
   assign soundFileAmplitudes [16041] = 8'd117;
   assign soundFileAmplitudes [16042] = 8'd119;
   assign soundFileAmplitudes [16043] = 8'd124;
   assign soundFileAmplitudes [16044] = 8'd127;
   assign soundFileAmplitudes [16045] = 8'd128;
   assign soundFileAmplitudes [16046] = 8'd128;
   assign soundFileAmplitudes [16047] = 8'd122;
   assign soundFileAmplitudes [16048] = 8'd122;
   assign soundFileAmplitudes [16049] = 8'd117;
   assign soundFileAmplitudes [16050] = 8'd112;
   assign soundFileAmplitudes [16051] = 8'd118;
   assign soundFileAmplitudes [16052] = 8'd121;
   assign soundFileAmplitudes [16053] = 8'd118;
   assign soundFileAmplitudes [16054] = 8'd126;
   assign soundFileAmplitudes [16055] = 8'd130;
   assign soundFileAmplitudes [16056] = 8'd133;
   assign soundFileAmplitudes [16057] = 8'd142;
   assign soundFileAmplitudes [16058] = 8'd143;
   assign soundFileAmplitudes [16059] = 8'd147;
   assign soundFileAmplitudes [16060] = 8'd146;
   assign soundFileAmplitudes [16061] = 8'd156;
   assign soundFileAmplitudes [16062] = 8'd158;
   assign soundFileAmplitudes [16063] = 8'd155;
   assign soundFileAmplitudes [16064] = 8'd140;
   assign soundFileAmplitudes [16065] = 8'd122;
   assign soundFileAmplitudes [16066] = 8'd120;
   assign soundFileAmplitudes [16067] = 8'd109;
   assign soundFileAmplitudes [16068] = 8'd101;
   assign soundFileAmplitudes [16069] = 8'd105;
   assign soundFileAmplitudes [16070] = 8'd107;
   assign soundFileAmplitudes [16071] = 8'd111;
   assign soundFileAmplitudes [16072] = 8'd112;
   assign soundFileAmplitudes [16073] = 8'd111;
   assign soundFileAmplitudes [16074] = 8'd123;
   assign soundFileAmplitudes [16075] = 8'd129;
   assign soundFileAmplitudes [16076] = 8'd144;
   assign soundFileAmplitudes [16077] = 8'd141;
   assign soundFileAmplitudes [16078] = 8'd128;
   assign soundFileAmplitudes [16079] = 8'd135;
   assign soundFileAmplitudes [16080] = 8'd142;
   assign soundFileAmplitudes [16081] = 8'd135;
   assign soundFileAmplitudes [16082] = 8'd114;
   assign soundFileAmplitudes [16083] = 8'd106;
   assign soundFileAmplitudes [16084] = 8'd113;
   assign soundFileAmplitudes [16085] = 8'd122;
   assign soundFileAmplitudes [16086] = 8'd120;
   assign soundFileAmplitudes [16087] = 8'd114;
   assign soundFileAmplitudes [16088] = 8'd101;
   assign soundFileAmplitudes [16089] = 8'd101;
   assign soundFileAmplitudes [16090] = 8'd117;
   assign soundFileAmplitudes [16091] = 8'd133;
   assign soundFileAmplitudes [16092] = 8'd141;
   assign soundFileAmplitudes [16093] = 8'd150;
   assign soundFileAmplitudes [16094] = 8'd153;
   assign soundFileAmplitudes [16095] = 8'd149;
   assign soundFileAmplitudes [16096] = 8'd145;
   assign soundFileAmplitudes [16097] = 8'd141;
   assign soundFileAmplitudes [16098] = 8'd140;
   assign soundFileAmplitudes [16099] = 8'd138;
   assign soundFileAmplitudes [16100] = 8'd128;
   assign soundFileAmplitudes [16101] = 8'd123;
   assign soundFileAmplitudes [16102] = 8'd108;
   assign soundFileAmplitudes [16103] = 8'd98;
   assign soundFileAmplitudes [16104] = 8'd112;
   assign soundFileAmplitudes [16105] = 8'd116;
   assign soundFileAmplitudes [16106] = 8'd117;
   assign soundFileAmplitudes [16107] = 8'd119;
   assign soundFileAmplitudes [16108] = 8'd120;
   assign soundFileAmplitudes [16109] = 8'd128;
   assign soundFileAmplitudes [16110] = 8'd126;
   assign soundFileAmplitudes [16111] = 8'd114;
   assign soundFileAmplitudes [16112] = 8'd122;
   assign soundFileAmplitudes [16113] = 8'd125;
   assign soundFileAmplitudes [16114] = 8'd133;
   assign soundFileAmplitudes [16115] = 8'd128;
   assign soundFileAmplitudes [16116] = 8'd119;
   assign soundFileAmplitudes [16117] = 8'd124;
   assign soundFileAmplitudes [16118] = 8'd127;
   assign soundFileAmplitudes [16119] = 8'd137;
   assign soundFileAmplitudes [16120] = 8'd132;
   assign soundFileAmplitudes [16121] = 8'd128;
   assign soundFileAmplitudes [16122] = 8'd126;
   assign soundFileAmplitudes [16123] = 8'd124;
   assign soundFileAmplitudes [16124] = 8'd121;
   assign soundFileAmplitudes [16125] = 8'd123;
   assign soundFileAmplitudes [16126] = 8'd127;
   assign soundFileAmplitudes [16127] = 8'd144;
   assign soundFileAmplitudes [16128] = 8'd148;
   assign soundFileAmplitudes [16129] = 8'd144;
   assign soundFileAmplitudes [16130] = 8'd140;
   assign soundFileAmplitudes [16131] = 8'd123;
   assign soundFileAmplitudes [16132] = 8'd118;
   assign soundFileAmplitudes [16133] = 8'd128;
   assign soundFileAmplitudes [16134] = 8'd128;
   assign soundFileAmplitudes [16135] = 8'd126;
   assign soundFileAmplitudes [16136] = 8'd130;
   assign soundFileAmplitudes [16137] = 8'd128;
   assign soundFileAmplitudes [16138] = 8'd121;
   assign soundFileAmplitudes [16139] = 8'd107;
   assign soundFileAmplitudes [16140] = 8'd112;
   assign soundFileAmplitudes [16141] = 8'd120;
   assign soundFileAmplitudes [16142] = 8'd127;
   assign soundFileAmplitudes [16143] = 8'd130;
   assign soundFileAmplitudes [16144] = 8'd120;
   assign soundFileAmplitudes [16145] = 8'd129;
   assign soundFileAmplitudes [16146] = 8'd122;
   assign soundFileAmplitudes [16147] = 8'd126;
   assign soundFileAmplitudes [16148] = 8'd127;
   assign soundFileAmplitudes [16149] = 8'd111;
   assign soundFileAmplitudes [16150] = 8'd131;
   assign soundFileAmplitudes [16151] = 8'd146;
   assign soundFileAmplitudes [16152] = 8'd143;
   assign soundFileAmplitudes [16153] = 8'd140;
   assign soundFileAmplitudes [16154] = 8'd133;
   assign soundFileAmplitudes [16155] = 8'd134;
   assign soundFileAmplitudes [16156] = 8'd141;
   assign soundFileAmplitudes [16157] = 8'd139;
   assign soundFileAmplitudes [16158] = 8'd141;
   assign soundFileAmplitudes [16159] = 8'd138;
   assign soundFileAmplitudes [16160] = 8'd129;
   assign soundFileAmplitudes [16161] = 8'd114;
   assign soundFileAmplitudes [16162] = 8'd111;
   assign soundFileAmplitudes [16163] = 8'd115;
   assign soundFileAmplitudes [16164] = 8'd115;
   assign soundFileAmplitudes [16165] = 8'd120;
   assign soundFileAmplitudes [16166] = 8'd115;
   assign soundFileAmplitudes [16167] = 8'd108;
   assign soundFileAmplitudes [16168] = 8'd115;
   assign soundFileAmplitudes [16169] = 8'd130;
   assign soundFileAmplitudes [16170] = 8'd139;
   assign soundFileAmplitudes [16171] = 8'd151;
   assign soundFileAmplitudes [16172] = 8'd146;
   assign soundFileAmplitudes [16173] = 8'd135;
   assign soundFileAmplitudes [16174] = 8'd117;
   assign soundFileAmplitudes [16175] = 8'd116;
   assign soundFileAmplitudes [16176] = 8'd123;
   assign soundFileAmplitudes [16177] = 8'd115;
   assign soundFileAmplitudes [16178] = 8'd123;
   assign soundFileAmplitudes [16179] = 8'd112;
   assign soundFileAmplitudes [16180] = 8'd111;
   assign soundFileAmplitudes [16181] = 8'd114;
   assign soundFileAmplitudes [16182] = 8'd107;
   assign soundFileAmplitudes [16183] = 8'd117;
   assign soundFileAmplitudes [16184] = 8'd128;
   assign soundFileAmplitudes [16185] = 8'd128;
   assign soundFileAmplitudes [16186] = 8'd136;
   assign soundFileAmplitudes [16187] = 8'd145;
   assign soundFileAmplitudes [16188] = 8'd141;
   assign soundFileAmplitudes [16189] = 8'd145;
   assign soundFileAmplitudes [16190] = 8'd145;
   assign soundFileAmplitudes [16191] = 8'd151;
   assign soundFileAmplitudes [16192] = 8'd155;
   assign soundFileAmplitudes [16193] = 8'd133;
   assign soundFileAmplitudes [16194] = 8'd123;
   assign soundFileAmplitudes [16195] = 8'd113;
   assign soundFileAmplitudes [16196] = 8'd108;
   assign soundFileAmplitudes [16197] = 8'd113;
   assign soundFileAmplitudes [16198] = 8'd100;
   assign soundFileAmplitudes [16199] = 8'd92;
   assign soundFileAmplitudes [16200] = 8'd94;
   assign soundFileAmplitudes [16201] = 8'd103;
   assign soundFileAmplitudes [16202] = 8'd113;
   assign soundFileAmplitudes [16203] = 8'd119;
   assign soundFileAmplitudes [16204] = 8'd133;
   assign soundFileAmplitudes [16205] = 8'd141;
   assign soundFileAmplitudes [16206] = 8'd135;
   assign soundFileAmplitudes [16207] = 8'd137;
   assign soundFileAmplitudes [16208] = 8'd144;
   assign soundFileAmplitudes [16209] = 8'd145;
   assign soundFileAmplitudes [16210] = 8'd140;
   assign soundFileAmplitudes [16211] = 8'd134;
   assign soundFileAmplitudes [16212] = 8'd128;
   assign soundFileAmplitudes [16213] = 8'd119;
   assign soundFileAmplitudes [16214] = 8'd111;
   assign soundFileAmplitudes [16215] = 8'd117;
   assign soundFileAmplitudes [16216] = 8'd133;
   assign soundFileAmplitudes [16217] = 8'd131;
   assign soundFileAmplitudes [16218] = 8'd124;
   assign soundFileAmplitudes [16219] = 8'd122;
   assign soundFileAmplitudes [16220] = 8'd127;
   assign soundFileAmplitudes [16221] = 8'd129;
   assign soundFileAmplitudes [16222] = 8'd142;
   assign soundFileAmplitudes [16223] = 8'd153;
   assign soundFileAmplitudes [16224] = 8'd154;
   assign soundFileAmplitudes [16225] = 8'd146;
   assign soundFileAmplitudes [16226] = 8'd129;
   assign soundFileAmplitudes [16227] = 8'd124;
   assign soundFileAmplitudes [16228] = 8'd128;
   assign soundFileAmplitudes [16229] = 8'd129;
   assign soundFileAmplitudes [16230] = 8'd117;
   assign soundFileAmplitudes [16231] = 8'd99;
   assign soundFileAmplitudes [16232] = 8'd75;
   assign soundFileAmplitudes [16233] = 8'd81;
   assign soundFileAmplitudes [16234] = 8'd102;
   assign soundFileAmplitudes [16235] = 8'd113;
   assign soundFileAmplitudes [16236] = 8'd118;
   assign soundFileAmplitudes [16237] = 8'd118;
   assign soundFileAmplitudes [16238] = 8'd111;
   assign soundFileAmplitudes [16239] = 8'd108;
   assign soundFileAmplitudes [16240] = 8'd138;
   assign soundFileAmplitudes [16241] = 8'd146;
   assign soundFileAmplitudes [16242] = 8'd157;
   assign soundFileAmplitudes [16243] = 8'd155;
   assign soundFileAmplitudes [16244] = 8'd146;
   assign soundFileAmplitudes [16245] = 8'd148;
   assign soundFileAmplitudes [16246] = 8'd127;
   assign soundFileAmplitudes [16247] = 8'd128;
   assign soundFileAmplitudes [16248] = 8'd141;
   assign soundFileAmplitudes [16249] = 8'd147;
   assign soundFileAmplitudes [16250] = 8'd134;
   assign soundFileAmplitudes [16251] = 8'd125;
   assign soundFileAmplitudes [16252] = 8'd122;
   assign soundFileAmplitudes [16253] = 8'd124;
   assign soundFileAmplitudes [16254] = 8'd126;
   assign soundFileAmplitudes [16255] = 8'd128;
   assign soundFileAmplitudes [16256] = 8'd140;
   assign soundFileAmplitudes [16257] = 8'd145;
   assign soundFileAmplitudes [16258] = 8'd145;
   assign soundFileAmplitudes [16259] = 8'd130;
   assign soundFileAmplitudes [16260] = 8'd123;
   assign soundFileAmplitudes [16261] = 8'd120;
   assign soundFileAmplitudes [16262] = 8'd123;
   assign soundFileAmplitudes [16263] = 8'd118;
   assign soundFileAmplitudes [16264] = 8'd111;
   assign soundFileAmplitudes [16265] = 8'd102;
   assign soundFileAmplitudes [16266] = 8'd102;
   assign soundFileAmplitudes [16267] = 8'd103;
   assign soundFileAmplitudes [16268] = 8'd112;
   assign soundFileAmplitudes [16269] = 8'd119;
   assign soundFileAmplitudes [16270] = 8'd115;
   assign soundFileAmplitudes [16271] = 8'd117;
   assign soundFileAmplitudes [16272] = 8'd118;
   assign soundFileAmplitudes [16273] = 8'd126;
   assign soundFileAmplitudes [16274] = 8'd123;
   assign soundFileAmplitudes [16275] = 8'd129;
   assign soundFileAmplitudes [16276] = 8'd126;
   assign soundFileAmplitudes [16277] = 8'd136;
   assign soundFileAmplitudes [16278] = 8'd143;
   assign soundFileAmplitudes [16279] = 8'd133;
   assign soundFileAmplitudes [16280] = 8'd148;
   assign soundFileAmplitudes [16281] = 8'd148;
   assign soundFileAmplitudes [16282] = 8'd137;
   assign soundFileAmplitudes [16283] = 8'd130;
   assign soundFileAmplitudes [16284] = 8'd135;
   assign soundFileAmplitudes [16285] = 8'd133;
   assign soundFileAmplitudes [16286] = 8'd135;
   assign soundFileAmplitudes [16287] = 8'd134;
   assign soundFileAmplitudes [16288] = 8'd127;
   assign soundFileAmplitudes [16289] = 8'd142;
   assign soundFileAmplitudes [16290] = 8'd136;
   assign soundFileAmplitudes [16291] = 8'd124;
   assign soundFileAmplitudes [16292] = 8'd122;
   assign soundFileAmplitudes [16293] = 8'd126;
   assign soundFileAmplitudes [16294] = 8'd136;
   assign soundFileAmplitudes [16295] = 8'd140;
   assign soundFileAmplitudes [16296] = 8'd129;
   assign soundFileAmplitudes [16297] = 8'd122;
   assign soundFileAmplitudes [16298] = 8'd117;
   assign soundFileAmplitudes [16299] = 8'd115;
   assign soundFileAmplitudes [16300] = 8'd121;
   assign soundFileAmplitudes [16301] = 8'd128;
   assign soundFileAmplitudes [16302] = 8'd120;
   assign soundFileAmplitudes [16303] = 8'd108;
   assign soundFileAmplitudes [16304] = 8'd103;
   assign soundFileAmplitudes [16305] = 8'd116;
   assign soundFileAmplitudes [16306] = 8'd118;
   assign soundFileAmplitudes [16307] = 8'd122;
   assign soundFileAmplitudes [16308] = 8'd126;
   assign soundFileAmplitudes [16309] = 8'd117;
   assign soundFileAmplitudes [16310] = 8'd122;
   assign soundFileAmplitudes [16311] = 8'd108;
   assign soundFileAmplitudes [16312] = 8'd121;
   assign soundFileAmplitudes [16313] = 8'd141;
   assign soundFileAmplitudes [16314] = 8'd143;
   assign soundFileAmplitudes [16315] = 8'd142;
   assign soundFileAmplitudes [16316] = 8'd141;
   assign soundFileAmplitudes [16317] = 8'd139;
   assign soundFileAmplitudes [16318] = 8'd126;
   assign soundFileAmplitudes [16319] = 8'd123;
   assign soundFileAmplitudes [16320] = 8'd123;
   assign soundFileAmplitudes [16321] = 8'd129;
   assign soundFileAmplitudes [16322] = 8'd139;
   assign soundFileAmplitudes [16323] = 8'd135;
   assign soundFileAmplitudes [16324] = 8'd124;
   assign soundFileAmplitudes [16325] = 8'd118;
   assign soundFileAmplitudes [16326] = 8'd118;
   assign soundFileAmplitudes [16327] = 8'd121;
   assign soundFileAmplitudes [16328] = 8'd119;
   assign soundFileAmplitudes [16329] = 8'd120;
   assign soundFileAmplitudes [16330] = 8'd125;
   assign soundFileAmplitudes [16331] = 8'd133;
   assign soundFileAmplitudes [16332] = 8'd131;
   assign soundFileAmplitudes [16333] = 8'd131;
   assign soundFileAmplitudes [16334] = 8'd128;
   assign soundFileAmplitudes [16335] = 8'd123;
   assign soundFileAmplitudes [16336] = 8'd121;
   assign soundFileAmplitudes [16337] = 8'd127;
   assign soundFileAmplitudes [16338] = 8'd127;
   assign soundFileAmplitudes [16339] = 8'd117;
   assign soundFileAmplitudes [16340] = 8'd121;
   assign soundFileAmplitudes [16341] = 8'd115;
   assign soundFileAmplitudes [16342] = 8'd121;
   assign soundFileAmplitudes [16343] = 8'd124;
   assign soundFileAmplitudes [16344] = 8'd121;
   assign soundFileAmplitudes [16345] = 8'd129;
   assign soundFileAmplitudes [16346] = 8'd128;
   assign soundFileAmplitudes [16347] = 8'd123;
   assign soundFileAmplitudes [16348] = 8'd132;
   assign soundFileAmplitudes [16349] = 8'd136;
   assign soundFileAmplitudes [16350] = 8'd134;
   assign soundFileAmplitudes [16351] = 8'd130;
   assign soundFileAmplitudes [16352] = 8'd130;
   assign soundFileAmplitudes [16353] = 8'd134;
   assign soundFileAmplitudes [16354] = 8'd130;
   assign soundFileAmplitudes [16355] = 8'd131;
   assign soundFileAmplitudes [16356] = 8'd120;
   assign soundFileAmplitudes [16357] = 8'd112;
   assign soundFileAmplitudes [16358] = 8'd118;
   assign soundFileAmplitudes [16359] = 8'd122;
   assign soundFileAmplitudes [16360] = 8'd125;
   assign soundFileAmplitudes [16361] = 8'd127;
   assign soundFileAmplitudes [16362] = 8'd114;
   assign soundFileAmplitudes [16363] = 8'd115;
   assign soundFileAmplitudes [16364] = 8'd120;
   assign soundFileAmplitudes [16365] = 8'd127;
   assign soundFileAmplitudes [16366] = 8'd142;
   assign soundFileAmplitudes [16367] = 8'd141;
   assign soundFileAmplitudes [16368] = 8'd130;
   assign soundFileAmplitudes [16369] = 8'd121;
   assign soundFileAmplitudes [16370] = 8'd129;
   assign soundFileAmplitudes [16371] = 8'd134;
   assign soundFileAmplitudes [16372] = 8'd137;
   assign soundFileAmplitudes [16373] = 8'd135;
   assign soundFileAmplitudes [16374] = 8'd119;
   assign soundFileAmplitudes [16375] = 8'd116;
   assign soundFileAmplitudes [16376] = 8'd112;
   assign soundFileAmplitudes [16377] = 8'd121;
   assign soundFileAmplitudes [16378] = 8'd139;
   assign soundFileAmplitudes [16379] = 8'd140;
   assign soundFileAmplitudes [16380] = 8'd129;
   assign soundFileAmplitudes [16381] = 8'd124;
   assign soundFileAmplitudes [16382] = 8'd122;
   assign soundFileAmplitudes [16383] = 8'd125;
   assign soundFileAmplitudes [16384] = 8'd139;
   assign soundFileAmplitudes [16385] = 8'd142;
   assign soundFileAmplitudes [16386] = 8'd134;
   assign soundFileAmplitudes [16387] = 8'd128;
   assign soundFileAmplitudes [16388] = 8'd126;
   assign soundFileAmplitudes [16389] = 8'd117;
   assign soundFileAmplitudes [16390] = 8'd115;
   assign soundFileAmplitudes [16391] = 8'd123;
   assign soundFileAmplitudes [16392] = 8'd125;
   assign soundFileAmplitudes [16393] = 8'd121;
   assign soundFileAmplitudes [16394] = 8'd111;
   assign soundFileAmplitudes [16395] = 8'd107;
   assign soundFileAmplitudes [16396] = 8'd111;
   assign soundFileAmplitudes [16397] = 8'd122;
   assign soundFileAmplitudes [16398] = 8'd129;
   assign soundFileAmplitudes [16399] = 8'd133;
   assign soundFileAmplitudes [16400] = 8'd130;
   assign soundFileAmplitudes [16401] = 8'd130;
   assign soundFileAmplitudes [16402] = 8'd131;
   assign soundFileAmplitudes [16403] = 8'd135;
   assign soundFileAmplitudes [16404] = 8'd140;
   assign soundFileAmplitudes [16405] = 8'd140;
   assign soundFileAmplitudes [16406] = 8'd140;
   assign soundFileAmplitudes [16407] = 8'd132;
   assign soundFileAmplitudes [16408] = 8'd133;
   assign soundFileAmplitudes [16409] = 8'd128;
   assign soundFileAmplitudes [16410] = 8'd124;
   assign soundFileAmplitudes [16411] = 8'd126;
   assign soundFileAmplitudes [16412] = 8'd124;
   assign soundFileAmplitudes [16413] = 8'd126;
   assign soundFileAmplitudes [16414] = 8'd133;
   assign soundFileAmplitudes [16415] = 8'd135;
   assign soundFileAmplitudes [16416] = 8'd135;
   assign soundFileAmplitudes [16417] = 8'd131;
   assign soundFileAmplitudes [16418] = 8'd123;
   assign soundFileAmplitudes [16419] = 8'd135;
   assign soundFileAmplitudes [16420] = 8'd145;
   assign soundFileAmplitudes [16421] = 8'd139;
   assign soundFileAmplitudes [16422] = 8'd123;
   assign soundFileAmplitudes [16423] = 8'd121;
   assign soundFileAmplitudes [16424] = 8'd115;
   assign soundFileAmplitudes [16425] = 8'd103;
   assign soundFileAmplitudes [16426] = 8'd103;
   assign soundFileAmplitudes [16427] = 8'd103;
   assign soundFileAmplitudes [16428] = 8'd105;
   assign soundFileAmplitudes [16429] = 8'd111;
   assign soundFileAmplitudes [16430] = 8'd115;
   assign soundFileAmplitudes [16431] = 8'd120;
   assign soundFileAmplitudes [16432] = 8'd127;
   assign soundFileAmplitudes [16433] = 8'd121;
   assign soundFileAmplitudes [16434] = 8'd123;
   assign soundFileAmplitudes [16435] = 8'd127;
   assign soundFileAmplitudes [16436] = 8'd143;
   assign soundFileAmplitudes [16437] = 8'd154;
   assign soundFileAmplitudes [16438] = 8'd157;
   assign soundFileAmplitudes [16439] = 8'd148;
   assign soundFileAmplitudes [16440] = 8'd131;
   assign soundFileAmplitudes [16441] = 8'd136;
   assign soundFileAmplitudes [16442] = 8'd133;
   assign soundFileAmplitudes [16443] = 8'd135;
   assign soundFileAmplitudes [16444] = 8'd133;
   assign soundFileAmplitudes [16445] = 8'd123;
   assign soundFileAmplitudes [16446] = 8'd113;
   assign soundFileAmplitudes [16447] = 8'd107;
   assign soundFileAmplitudes [16448] = 8'd113;
   assign soundFileAmplitudes [16449] = 8'd125;
   assign soundFileAmplitudes [16450] = 8'd132;
   assign soundFileAmplitudes [16451] = 8'd130;
   assign soundFileAmplitudes [16452] = 8'd129;
   assign soundFileAmplitudes [16453] = 8'd118;
   assign soundFileAmplitudes [16454] = 8'd121;
   assign soundFileAmplitudes [16455] = 8'd132;
   assign soundFileAmplitudes [16456] = 8'd140;
   assign soundFileAmplitudes [16457] = 8'd136;
   assign soundFileAmplitudes [16458] = 8'd128;
   assign soundFileAmplitudes [16459] = 8'd124;
   assign soundFileAmplitudes [16460] = 8'd112;
   assign soundFileAmplitudes [16461] = 8'd104;
   assign soundFileAmplitudes [16462] = 8'd108;
   assign soundFileAmplitudes [16463] = 8'd111;
   assign soundFileAmplitudes [16464] = 8'd115;
   assign soundFileAmplitudes [16465] = 8'd119;
   assign soundFileAmplitudes [16466] = 8'd110;
   assign soundFileAmplitudes [16467] = 8'd118;
   assign soundFileAmplitudes [16468] = 8'd119;
   assign soundFileAmplitudes [16469] = 8'd127;
   assign soundFileAmplitudes [16470] = 8'd137;
   assign soundFileAmplitudes [16471] = 8'd137;
   assign soundFileAmplitudes [16472] = 8'd149;
   assign soundFileAmplitudes [16473] = 8'd152;
   assign soundFileAmplitudes [16474] = 8'd151;
   assign soundFileAmplitudes [16475] = 8'd149;
   assign soundFileAmplitudes [16476] = 8'd142;
   assign soundFileAmplitudes [16477] = 8'd134;
   assign soundFileAmplitudes [16478] = 8'd135;
   assign soundFileAmplitudes [16479] = 8'd123;
   assign soundFileAmplitudes [16480] = 8'd115;
   assign soundFileAmplitudes [16481] = 8'd115;
   assign soundFileAmplitudes [16482] = 8'd109;
   assign soundFileAmplitudes [16483] = 8'd114;
   assign soundFileAmplitudes [16484] = 8'd117;
   assign soundFileAmplitudes [16485] = 8'd114;
   assign soundFileAmplitudes [16486] = 8'd115;
   assign soundFileAmplitudes [16487] = 8'd119;
   assign soundFileAmplitudes [16488] = 8'd121;
   assign soundFileAmplitudes [16489] = 8'd128;
   assign soundFileAmplitudes [16490] = 8'd138;
   assign soundFileAmplitudes [16491] = 8'd138;
   assign soundFileAmplitudes [16492] = 8'd131;
   assign soundFileAmplitudes [16493] = 8'd124;
   assign soundFileAmplitudes [16494] = 8'd121;
   assign soundFileAmplitudes [16495] = 8'd113;
   assign soundFileAmplitudes [16496] = 8'd112;
   assign soundFileAmplitudes [16497] = 8'd115;
   assign soundFileAmplitudes [16498] = 8'd115;
   assign soundFileAmplitudes [16499] = 8'd116;
   assign soundFileAmplitudes [16500] = 8'd115;
   assign soundFileAmplitudes [16501] = 8'd107;
   assign soundFileAmplitudes [16502] = 8'd118;
   assign soundFileAmplitudes [16503] = 8'd134;
   assign soundFileAmplitudes [16504] = 8'd138;
   assign soundFileAmplitudes [16505] = 8'd139;
   assign soundFileAmplitudes [16506] = 8'd140;
   assign soundFileAmplitudes [16507] = 8'd145;
   assign soundFileAmplitudes [16508] = 8'd155;
   assign soundFileAmplitudes [16509] = 8'd161;
   assign soundFileAmplitudes [16510] = 8'd145;
   assign soundFileAmplitudes [16511] = 8'd144;
   assign soundFileAmplitudes [16512] = 8'd142;
   assign soundFileAmplitudes [16513] = 8'd136;
   assign soundFileAmplitudes [16514] = 8'd129;
   assign soundFileAmplitudes [16515] = 8'd116;
   assign soundFileAmplitudes [16516] = 8'd109;
   assign soundFileAmplitudes [16517] = 8'd105;
   assign soundFileAmplitudes [16518] = 8'd106;
   assign soundFileAmplitudes [16519] = 8'd109;
   assign soundFileAmplitudes [16520] = 8'd119;
   assign soundFileAmplitudes [16521] = 8'd123;
   assign soundFileAmplitudes [16522] = 8'd121;
   assign soundFileAmplitudes [16523] = 8'd113;
   assign soundFileAmplitudes [16524] = 8'd125;
   assign soundFileAmplitudes [16525] = 8'd138;
   assign soundFileAmplitudes [16526] = 8'd143;
   assign soundFileAmplitudes [16527] = 8'd133;
   assign soundFileAmplitudes [16528] = 8'd128;
   assign soundFileAmplitudes [16529] = 8'd129;
   assign soundFileAmplitudes [16530] = 8'd114;
   assign soundFileAmplitudes [16531] = 8'd115;
   assign soundFileAmplitudes [16532] = 8'd117;
   assign soundFileAmplitudes [16533] = 8'd117;
   assign soundFileAmplitudes [16534] = 8'd119;
   assign soundFileAmplitudes [16535] = 8'd121;
   assign soundFileAmplitudes [16536] = 8'd116;
   assign soundFileAmplitudes [16537] = 8'd113;
   assign soundFileAmplitudes [16538] = 8'd118;
   assign soundFileAmplitudes [16539] = 8'd128;
   assign soundFileAmplitudes [16540] = 8'd144;
   assign soundFileAmplitudes [16541] = 8'd146;
   assign soundFileAmplitudes [16542] = 8'd147;
   assign soundFileAmplitudes [16543] = 8'd153;
   assign soundFileAmplitudes [16544] = 8'd146;
   assign soundFileAmplitudes [16545] = 8'd145;
   assign soundFileAmplitudes [16546] = 8'd151;
   assign soundFileAmplitudes [16547] = 8'd149;
   assign soundFileAmplitudes [16548] = 8'd142;
   assign soundFileAmplitudes [16549] = 8'd132;
   assign soundFileAmplitudes [16550] = 8'd114;
   assign soundFileAmplitudes [16551] = 8'd97;
   assign soundFileAmplitudes [16552] = 8'd94;
   assign soundFileAmplitudes [16553] = 8'd100;
   assign soundFileAmplitudes [16554] = 8'd119;
   assign soundFileAmplitudes [16555] = 8'd128;
   assign soundFileAmplitudes [16556] = 8'd125;
   assign soundFileAmplitudes [16557] = 8'd116;
   assign soundFileAmplitudes [16558] = 8'd120;
   assign soundFileAmplitudes [16559] = 8'd137;
   assign soundFileAmplitudes [16560] = 8'd143;
   assign soundFileAmplitudes [16561] = 8'd147;
   assign soundFileAmplitudes [16562] = 8'd139;
   assign soundFileAmplitudes [16563] = 8'd134;
   assign soundFileAmplitudes [16564] = 8'd121;
   assign soundFileAmplitudes [16565] = 8'd110;
   assign soundFileAmplitudes [16566] = 8'd119;
   assign soundFileAmplitudes [16567] = 8'd129;
   assign soundFileAmplitudes [16568] = 8'd126;
   assign soundFileAmplitudes [16569] = 8'd115;
   assign soundFileAmplitudes [16570] = 8'd108;
   assign soundFileAmplitudes [16571] = 8'd113;
   assign soundFileAmplitudes [16572] = 8'd125;
   assign soundFileAmplitudes [16573] = 8'd125;
   assign soundFileAmplitudes [16574] = 8'd130;
   assign soundFileAmplitudes [16575] = 8'd123;
   assign soundFileAmplitudes [16576] = 8'd123;
   assign soundFileAmplitudes [16577] = 8'd141;
   assign soundFileAmplitudes [16578] = 8'd142;
   assign soundFileAmplitudes [16579] = 8'd141;
   assign soundFileAmplitudes [16580] = 8'd144;
   assign soundFileAmplitudes [16581] = 8'd143;
   assign soundFileAmplitudes [16582] = 8'd135;
   assign soundFileAmplitudes [16583] = 8'd130;
   assign soundFileAmplitudes [16584] = 8'd122;
   assign soundFileAmplitudes [16585] = 8'd111;
   assign soundFileAmplitudes [16586] = 8'd110;
   assign soundFileAmplitudes [16587] = 8'd106;
   assign soundFileAmplitudes [16588] = 8'd119;
   assign soundFileAmplitudes [16589] = 8'd126;
   assign soundFileAmplitudes [16590] = 8'd122;
   assign soundFileAmplitudes [16591] = 8'd117;
   assign soundFileAmplitudes [16592] = 8'd120;
   assign soundFileAmplitudes [16593] = 8'd145;
   assign soundFileAmplitudes [16594] = 8'd154;
   assign soundFileAmplitudes [16595] = 8'd150;
   assign soundFileAmplitudes [16596] = 8'd135;
   assign soundFileAmplitudes [16597] = 8'd125;
   assign soundFileAmplitudes [16598] = 8'd116;
   assign soundFileAmplitudes [16599] = 8'd110;
   assign soundFileAmplitudes [16600] = 8'd115;
   assign soundFileAmplitudes [16601] = 8'd121;
   assign soundFileAmplitudes [16602] = 8'd123;
   assign soundFileAmplitudes [16603] = 8'd124;
   assign soundFileAmplitudes [16604] = 8'd120;
   assign soundFileAmplitudes [16605] = 8'd120;
   assign soundFileAmplitudes [16606] = 8'd127;
   assign soundFileAmplitudes [16607] = 8'd134;
   assign soundFileAmplitudes [16608] = 8'd140;
   assign soundFileAmplitudes [16609] = 8'd137;
   assign soundFileAmplitudes [16610] = 8'd131;
   assign soundFileAmplitudes [16611] = 8'd128;
   assign soundFileAmplitudes [16612] = 8'd136;
   assign soundFileAmplitudes [16613] = 8'd132;
   assign soundFileAmplitudes [16614] = 8'd130;
   assign soundFileAmplitudes [16615] = 8'd132;
   assign soundFileAmplitudes [16616] = 8'd130;
   assign soundFileAmplitudes [16617] = 8'd123;
   assign soundFileAmplitudes [16618] = 8'd113;
   assign soundFileAmplitudes [16619] = 8'd103;
   assign soundFileAmplitudes [16620] = 8'd99;
   assign soundFileAmplitudes [16621] = 8'd106;
   assign soundFileAmplitudes [16622] = 8'd116;
   assign soundFileAmplitudes [16623] = 8'd125;
   assign soundFileAmplitudes [16624] = 8'd124;
   assign soundFileAmplitudes [16625] = 8'd124;
   assign soundFileAmplitudes [16626] = 8'd118;
   assign soundFileAmplitudes [16627] = 8'd123;
   assign soundFileAmplitudes [16628] = 8'd144;
   assign soundFileAmplitudes [16629] = 8'd148;
   assign soundFileAmplitudes [16630] = 8'd135;
   assign soundFileAmplitudes [16631] = 8'd132;
   assign soundFileAmplitudes [16632] = 8'd126;
   assign soundFileAmplitudes [16633] = 8'd110;
   assign soundFileAmplitudes [16634] = 8'd113;
   assign soundFileAmplitudes [16635] = 8'd122;
   assign soundFileAmplitudes [16636] = 8'd129;
   assign soundFileAmplitudes [16637] = 8'd133;
   assign soundFileAmplitudes [16638] = 8'd135;
   assign soundFileAmplitudes [16639] = 8'd127;
   assign soundFileAmplitudes [16640] = 8'd130;
   assign soundFileAmplitudes [16641] = 8'd136;
   assign soundFileAmplitudes [16642] = 8'd137;
   assign soundFileAmplitudes [16643] = 8'd143;
   assign soundFileAmplitudes [16644] = 8'd138;
   assign soundFileAmplitudes [16645] = 8'd133;
   assign soundFileAmplitudes [16646] = 8'd135;
   assign soundFileAmplitudes [16647] = 8'd142;
   assign soundFileAmplitudes [16648] = 8'd123;
   assign soundFileAmplitudes [16649] = 8'd114;
   assign soundFileAmplitudes [16650] = 8'd119;
   assign soundFileAmplitudes [16651] = 8'd125;
   assign soundFileAmplitudes [16652] = 8'd124;
   assign soundFileAmplitudes [16653] = 8'd114;
   assign soundFileAmplitudes [16654] = 8'd108;
   assign soundFileAmplitudes [16655] = 8'd103;
   assign soundFileAmplitudes [16656] = 8'd115;
   assign soundFileAmplitudes [16657] = 8'd129;
   assign soundFileAmplitudes [16658] = 8'd132;
   assign soundFileAmplitudes [16659] = 8'd132;
   assign soundFileAmplitudes [16660] = 8'd124;
   assign soundFileAmplitudes [16661] = 8'd121;
   assign soundFileAmplitudes [16662] = 8'd139;
   assign soundFileAmplitudes [16663] = 8'd147;
   assign soundFileAmplitudes [16664] = 8'd136;
   assign soundFileAmplitudes [16665] = 8'd121;
   assign soundFileAmplitudes [16666] = 8'd122;
   assign soundFileAmplitudes [16667] = 8'd116;
   assign soundFileAmplitudes [16668] = 8'd110;
   assign soundFileAmplitudes [16669] = 8'd119;
   assign soundFileAmplitudes [16670] = 8'd122;
   assign soundFileAmplitudes [16671] = 8'd125;
   assign soundFileAmplitudes [16672] = 8'd135;
   assign soundFileAmplitudes [16673] = 8'd132;
   assign soundFileAmplitudes [16674] = 8'd130;
   assign soundFileAmplitudes [16675] = 8'd139;
   assign soundFileAmplitudes [16676] = 8'd136;
   assign soundFileAmplitudes [16677] = 8'd144;
   assign soundFileAmplitudes [16678] = 8'd140;
   assign soundFileAmplitudes [16679] = 8'd139;
   assign soundFileAmplitudes [16680] = 8'd140;
   assign soundFileAmplitudes [16681] = 8'd136;
   assign soundFileAmplitudes [16682] = 8'd142;
   assign soundFileAmplitudes [16683] = 8'd128;
   assign soundFileAmplitudes [16684] = 8'd124;
   assign soundFileAmplitudes [16685] = 8'd124;
   assign soundFileAmplitudes [16686] = 8'd118;
   assign soundFileAmplitudes [16687] = 8'd112;
   assign soundFileAmplitudes [16688] = 8'd110;
   assign soundFileAmplitudes [16689] = 8'd105;
   assign soundFileAmplitudes [16690] = 8'd114;
   assign soundFileAmplitudes [16691] = 8'd131;
   assign soundFileAmplitudes [16692] = 8'd124;
   assign soundFileAmplitudes [16693] = 8'd125;
   assign soundFileAmplitudes [16694] = 8'd119;
   assign soundFileAmplitudes [16695] = 8'd125;
   assign soundFileAmplitudes [16696] = 8'd143;
   assign soundFileAmplitudes [16697] = 8'd154;
   assign soundFileAmplitudes [16698] = 8'd151;
   assign soundFileAmplitudes [16699] = 8'd135;
   assign soundFileAmplitudes [16700] = 8'd123;
   assign soundFileAmplitudes [16701] = 8'd110;
   assign soundFileAmplitudes [16702] = 8'd104;
   assign soundFileAmplitudes [16703] = 8'd110;
   assign soundFileAmplitudes [16704] = 8'd115;
   assign soundFileAmplitudes [16705] = 8'd120;
   assign soundFileAmplitudes [16706] = 8'd130;
   assign soundFileAmplitudes [16707] = 8'd123;
   assign soundFileAmplitudes [16708] = 8'd118;
   assign soundFileAmplitudes [16709] = 8'd120;
   assign soundFileAmplitudes [16710] = 8'd118;
   assign soundFileAmplitudes [16711] = 8'd129;
   assign soundFileAmplitudes [16712] = 8'd142;
   assign soundFileAmplitudes [16713] = 8'd149;
   assign soundFileAmplitudes [16714] = 8'd151;
   assign soundFileAmplitudes [16715] = 8'd143;
   assign soundFileAmplitudes [16716] = 8'd143;
   assign soundFileAmplitudes [16717] = 8'd142;
   assign soundFileAmplitudes [16718] = 8'd130;
   assign soundFileAmplitudes [16719] = 8'd123;
   assign soundFileAmplitudes [16720] = 8'd122;
   assign soundFileAmplitudes [16721] = 8'd118;
   assign soundFileAmplitudes [16722] = 8'd107;
   assign soundFileAmplitudes [16723] = 8'd83;
   assign soundFileAmplitudes [16724] = 8'd78;
   assign soundFileAmplitudes [16725] = 8'd104;
   assign soundFileAmplitudes [16726] = 8'd121;
   assign soundFileAmplitudes [16727] = 8'd129;
   assign soundFileAmplitudes [16728] = 8'd132;
   assign soundFileAmplitudes [16729] = 8'd131;
   assign soundFileAmplitudes [16730] = 8'd138;
   assign soundFileAmplitudes [16731] = 8'd156;
   assign soundFileAmplitudes [16732] = 8'd162;
   assign soundFileAmplitudes [16733] = 8'd145;
   assign soundFileAmplitudes [16734] = 8'd136;
   assign soundFileAmplitudes [16735] = 8'd134;
   assign soundFileAmplitudes [16736] = 8'd119;
   assign soundFileAmplitudes [16737] = 8'd109;
   assign soundFileAmplitudes [16738] = 8'd105;
   assign soundFileAmplitudes [16739] = 8'd105;
   assign soundFileAmplitudes [16740] = 8'd109;
   assign soundFileAmplitudes [16741] = 8'd119;
   assign soundFileAmplitudes [16742] = 8'd123;
   assign soundFileAmplitudes [16743] = 8'd132;
   assign soundFileAmplitudes [16744] = 8'd132;
   assign soundFileAmplitudes [16745] = 8'd132;
   assign soundFileAmplitudes [16746] = 8'd137;
   assign soundFileAmplitudes [16747] = 8'd150;
   assign soundFileAmplitudes [16748] = 8'd161;
endmodule
